----------------------------------------------------------------------------------
-- Engineer: Jozsef Laszlo ( rbendr AT gmail DOT com )
-- 
-- Create Date:    08:47:30 03/05/2017 
-- Design Name: 	 TVC Extra rom 
-- Module Name:    soundctrl - Behavioral 
-- Project Name:   TVC Home computer VHDL version
-- Description: 
--						 TVC Sound generator 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: All rights reserved
-- Status: works
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity extrom8k is
    Port ( CLK : in  STD_LOGIC;
             A : in  STD_LOGIC_VECTOR (12 downto 0);
          DOUT : out STD_LOGIC_VECTOR (7 downto 0)
		   );
				
end extrom8k;

architecture Behavioral of extrom8k is

type  
  romarray is array(0 to 8191) of std_logic_vector(7 downto 0);

constant
  myROM : romarray := (
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3E",x"D0",x"D3",x"02",x"3A",x"21",
x"0B",x"B7",x"20",x"04",x"08",x"32",x"1B",x"0B",x"21",x"6B",x"FB",x"11",x"40",x"07",
x"01",x"40",x"01",x"ED",x"B0",x"3E",x"40",x"E5",x"0E",x"0A",x"ED",x"B0",x"E1",x"3D",
x"20",x"F7",x"21",x"0E",x"FB",x"11",x"00",x"0B",x"0E",x"10",x"ED",x"B0",x"11",x"30",
x"00",x"0E",x"10",x"ED",x"B0",x"11",x"23",x"0B",x"0E",x"26",x"ED",x"B0",x"3E",x"FC",
x"32",x"10",x"0B",x"3E",x"80",x"32",x"13",x"0B",x"07",x"32",x"1F",x"0B",x"21",x"10",
x"0F",x"22",x"17",x"0B",x"DB",x"5A",x"01",x"03",x"04",x"21",x"40",x"00",x"57",x"3E",
x"04",x"90",x"0F",x"0F",x"D3",x"03",x"7A",x"A1",x"FE",x"03",x"E5",x"D9",x"28",x"11",
x"21",x"5C",x"FB",x"B7",x"28",x"1B",x"21",x"58",x"FB",x"3D",x"28",x"15",x"21",x"62",
x"FB",x"18",x"10",x"21",x"00",x"C0",x"11",x"54",x"FB",x"06",x"04",x"1A",x"BE",x"20",
x"0D",x"13",x"23",x"10",x"F8",x"4E",x"0C",x"06",x"00",x"D1",x"ED",x"B0",x"18",x"03",
x"E1",x"36",x"FF",x"D9",x"7A",x"0F",x"0F",x"11",x"30",x"00",x"19",x"10",x"B9",x"06",
x"04",x"57",x"A1",x"20",x"0B",x"3E",x"04",x"90",x"32",x"07",x"0B",x"32",x"0F",x"0B",
x"18",x"07",x"7A",x"0F",x"0F",x"10",x"EC",x"3E",x"FF",x"32",x"1C",x"0B",x"21",x"47",
x"00",x"11",x"30",x"00",x"06",x"04",x"AF",x"77",x"19",x"10",x"FC",x"1E",x"40",x"21",
x"70",x"00",x"D5",x"DD",x"E1",x"E5",x"FD",x"E1",x"46",x"04",x"1A",x"BE",x"20",x"07",
x"23",x"13",x"10",x"F8",x"FD",x"34",x"07",x"FD",x"E5",x"E1",x"11",x"30",x"00",x"19",
x"CB",x"44",x"28",x"0C",x"DD",x"E5",x"E1",x"19",x"CB",x"44",x"20",x"09",x"E5",x"DD",
x"E1",x"19",x"DD",x"E5",x"D1",x"18",x"D4",x"3E",x"F0",x"D3",x"02",x"CD",x"E8",x"FF",
x"DD",x"21",x"40",x"00",x"06",x"04",x"DB",x"5A",x"4F",x"3E",x"04",x"90",x"0F",x"0F",
x"D3",x"03",x"DD",x"7E",x"00",x"3C",x"28",x"15",x"79",x"E6",x"03",x"28",x"10",x"2A",
x"0B",x"C0",x"C5",x"DD",x"E5",x"CD",x"F9",x"FF",x"DD",x"E1",x"C1",x"3E",x"F0",x"D3",
x"02",x"11",x"30",x"00",x"DD",x"19",x"79",x"0F",x"0F",x"10",x"D3",x"21",x"D3",x"C2",
x"C3",x"F0",x"FF",x"08",x"3E",x"D0",x"D3",x"02",x"11",x"2E",x"FB",x"21",x"23",x"0B",
x"01",x"1E",x"00",x"1A",x"13",x"ED",x"A1",x"20",x"0B",x"EA",x"4B",x"F1",x"3A",x"21",
x"0B",x"B7",x"3E",x"FF",x"28",x"01",x"AF",x"32",x"21",x"0B",x"08",x"D3",x"02",x"C3",
x"3A",x"02",x"68",x"26",x"00",x"19",x"18",x"05",x"21",x"07",x"00",x"19",x"7E",x"FE",
x"04",x"30",x"64",x"D9",x"21",x"40",x"00",x"11",x"30",x"00",x"47",x"0F",x"0F",x"32",
x"11",x"0B",x"D3",x"03",x"78",x"B7",x"28",x"03",x"19",x"10",x"FD",x"7E",x"3C",x"28",
x"49",x"4E",x"23",x"11",x"5D",x"FB",x"1A",x"13",x"ED",x"A1",x"20",x"09",x"EA",x"94",
x"F1",x"D9",x"21",x"91",x"F2",x"18",x"04",x"D9",x"21",x"0D",x"C0",x"7E",x"3D",x"B9",
x"38",x"34",x"23",x"EB",x"69",x"26",x"00",x"29",x"19",x"5E",x"23",x"56",x"EB",x"3A",
x"11",x"0B",x"07",x"07",x"E6",x"03",x"DD",x"21",x"48",x"00",x"11",x"30",x"00",x"28",
x"05",x"47",x"DD",x"19",x"10",x"FC",x"08",x"D1",x"C1",x"CD",x"F9",x"FF",x"21",x"FC",
x"C3",x"C3",x"F0",x"FF",x"D9",x"3A",x"1C",x"0B",x"77",x"3E",x"FE",x"11",x"3E",x"FF",
x"D1",x"C1",x"18",x"EC",x"07",x"21",x"00",x"0B",x"11",x"0E",x"FB",x"DD",x"21",x"07",
x"0B",x"38",x"0A",x"21",x"08",x"0B",x"11",x"16",x"FB",x"DD",x"21",x"0F",x"0B",x"07",
x"07",x"07",x"E6",x"07",x"FE",x"07",x"28",x"12",x"4F",x"06",x"00",x"09",x"EB",x"09",
x"EB",x"7E",x"FE",x"06",x"CC",x"1E",x"F2",x"07",x"38",x"02",x"1A",x"77",x"21",x"0E",
x"C4",x"C3",x"F0",x"FF",x"08",x"3A",x"1C",x"0B",x"DD",x"77",x"00",x"08",x"C9",x"06",
x"04",x"CB",x"19",x"38",x"13",x"C5",x"3E",x"04",x"90",x"0F",x"0F",x"D3",x"03",x"2A",
x"0E",x"C0",x"CD",x"F9",x"FF",x"3E",x"F0",x"D3",x"02",x"C1",x"10",x"E7",x"3A",x"11",
x"0B",x"D3",x"03",x"E1",x"C3",x"F0",x"FF",x"EB",x"E5",x"D5",x"C5",x"E5",x"D5",x"EB",
x"2A",x"19",x"0B",x"B7",x"ED",x"52",x"3E",x"FA",x"D1",x"E1",x"D8",x"4E",x"EB",x"CD",
x"F9",x"FF",x"C1",x"D1",x"E1",x"B7",x"C0",x"ED",x"A1",x"E0",x"18",x"E0",x"E5",x"D5",
x"C5",x"E5",x"D5",x"2A",x"19",x"0B",x"B7",x"ED",x"52",x"3E",x"FA",x"D1",x"E1",x"D8",
x"CD",x"F9",x"FF",x"08",x"79",x"C1",x"D1",x"E1",x"08",x"B7",x"C0",x"08",x"12",x"AF",
x"EB",x"ED",x"A1",x"EB",x"E0",x"18",x"DB",x"05",x"05",x"F3",x"39",x"F3",x"B7",x"F3",
x"A4",x"F2",x"57",x"F3",x"32",x"69",x"0B",x"3E",x"EE",x"32",x"6A",x"0B",x"C5",x"E5",
x"3A",x"13",x"0B",x"E6",x"C3",x"32",x"13",x"0B",x"D3",x"06",x"3A",x"69",x"0B",x"FE",
x"09",x"38",x"02",x"3E",x"08",x"6F",x"26",x"00",x"29",x"11",x"C6",x"F3",x"19",x"5E",
x"23",x"56",x"7A",x"E6",x"0F",x"F6",x"10",x"57",x"3A",x"12",x"0B",x"E6",x"C0",x"B2",
x"32",x"12",x"0B",x"D3",x"05",x"7B",x"D3",x"04",x"3A",x"6A",x"0B",x"E6",x"B4",x"F6",
x"4A",x"67",x"01",x"11",x"04",x"11",x"03",x"40",x"DB",x"5A",x"6F",x"A3",x"20",x"0A",
x"ED",x"79",x"ED",x"79",x"ED",x"79",x"ED",x"51",x"ED",x"61",x"3E",x"10",x"81",x"4F",
x"7D",x"0F",x"0F",x"10",x"E9",x"AF",x"32",x"71",x"0B",x"E1",x"C1",x"C9",x"CD",x"31",
x"F3",x"C0",x"3A",x"14",x"0B",x"B7",x"20",x"F6",x"61",x"3A",x"11",x"0B",x"0F",x"0F",
x"E6",x"30",x"C6",x"11",x"4F",x"AF",x"3F",x"C9",x"00",x"CD",x"0A",x"F3",x"C0",x"ED",
x"78",x"E6",x"81",x"FE",x"81",x"3F",x"D8",x"CD",x"31",x"F3",x"28",x"F3",x"C9",x"3A",
x"16",x"0B",x"B7",x"C8",x"3E",x"F5",x"C9",x"FA",x"59",x"F3",x"CD",x"1F",x"F3",x"D0",
x"3A",x"71",x"0B",x"B7",x"C4",x"A4",x"F2",x"3E",x"05",x"ED",x"79",x"CD",x"31",x"F3",
x"C0",x"ED",x"78",x"0F",x"30",x"F7",x"0D",x"ED",x"61",x"AF",x"C9",x"CD",x"0A",x"F3",
x"D0",x"3A",x"71",x"0B",x"B7",x"C4",x"A4",x"F2",x"ED",x"78",x"0F",x"0F",x"30",x"06",
x"0D",x"ED",x"78",x"4F",x"AF",x"C9",x"F3",x"3A",x"11",x"0B",x"E6",x"F0",x"F6",x"07",
x"D3",x"03",x"3E",x"25",x"ED",x"79",x"DB",x"58",x"E6",x"18",x"20",x"09",x"21",x"62",
x"0B",x"CB",x"DE",x"3E",x"F5",x"FB",x"C9",x"ED",x"78",x"0F",x"0F",x"30",x"EB",x"3E",
x"05",x"ED",x"79",x"ED",x"78",x"0D",x"ED",x"60",x"FB",x"E6",x"38",x"28",x"14",x"47",
x"0C",x"3E",x"11",x"ED",x"79",x"3E",x"F4",x"CB",x"58",x"20",x"08",x"3E",x"F2",x"CB",
x"60",x"20",x"02",x"3E",x"F3",x"4C",x"C9",x"FA",x"C0",x"F3",x"21",x"3C",x"F3",x"C3",
x"4B",x"F2",x"21",x"59",x"F3",x"C3",x"6C",x"F2",x"88",x"0C",x"75",x"0D",x"BA",x"0E",
x"5D",x"0F",x"AF",x"0F",x"D7",x"0F",x"EC",x"0F",x"F6",x"0F",x"FB",x"0F",x"CD",x"93",
x"F5",x"18",x"17",x"CD",x"30",x"F6",x"18",x"12",x"CD",x"FA",x"F3",x"18",x"0D",x"CD",
x"58",x"F5",x"18",x"08",x"CD",x"05",x"F6",x"18",x"03",x"CD",x"07",x"F7",x"21",x"E7",
x"D9",x"C3",x"F0",x"FF",x"F2",x"CF",x"F4",x"CD",x"62",x"F7",x"3E",x"EB",x"C0",x"21",
x"F3",x"0B",x"01",x"21",x"01",x"CD",x"4F",x"F5",x"21",x"F4",x"0B",x"CD",x"26",x"F5",
x"CD",x"3C",x"F7",x"21",x"4E",x"F7",x"CD",x"30",x"F7",x"CD",x"3C",x"F7",x"3E",x"FF",
x"32",x"13",x"0D",x"21",x"05",x"0C",x"22",x"10",x"0D",x"21",x"00",x"01",x"22",x"09",
x"0D",x"AF",x"32",x"0B",x"0D",x"32",x"0C",x"0D",x"32",x"0D",x"0D",x"CD",x"7B",x"F7",
x"38",x"13",x"3A",x"0B",x"0D",x"FE",x"F5",x"20",x"D9",x"21",x"00",x"00",x"22",x"6F",
x"0B",x"21",x"F3",x"0B",x"36",x"00",x"C9",x"21",x"58",x"F7",x"D9",x"21",x"05",x"0C",
x"E5",x"11",x"F4",x"0B",x"1A",x"B7",x"28",x"0A",x"47",x"04",x"1A",x"96",x"20",x"08",
x"13",x"23",x"10",x"F8",x"21",x"44",x"F7",x"D9",x"D9",x"08",x"CD",x"30",x"F7",x"E1",
x"E5",x"7E",x"B7",x"C4",x"30",x"F7",x"CD",x"3C",x"F7",x"08",x"E1",x"20",x"9D",x"3A",
x"14",x"0D",x"B7",x"28",x"0E",x"21",x"0C",x"0D",x"7E",x"B7",x"28",x"07",x"AF",x"77",
x"3E",x"E6",x"C3",x"45",x"F4",x"3A",x"F3",x"0B",x"D6",x"11",x"32",x"6B",x"0B",x"3E",
x"00",x"32",x"13",x"0D",x"21",x"05",x"0C",x"11",x"F4",x"0B",x"7E",x"FE",x"11",x"38",
x"02",x"3E",x"10",x"3C",x"4F",x"06",x"00",x"ED",x"B0",x"21",x"05",x"0C",x"5E",x"1C",
x"16",x"00",x"19",x"22",x"07",x"0D",x"2A",x"05",x"0D",x"AF",x"ED",x"52",x"22",x"05",
x"0D",x"11",x"F4",x"0B",x"C3",x"B5",x"F5",x"CD",x"6B",x"F7",x"3E",x"EB",x"C0",x"3A",
x"0C",x"0D",x"B7",x"3E",x"E6",x"C0",x"21",x"14",x"0D",x"01",x"20",x"01",x"CD",x"4F",
x"F5",x"21",x"15",x"0D",x"CD",x"26",x"F5",x"3A",x"6B",x"0B",x"B7",x"3E",x"01",x"20",
x"02",x"3E",x"11",x"32",x"14",x"0D",x"32",x"2F",x"0E",x"21",x"6D",x"0B",x"7E",x"36",
x"00",x"32",x"30",x"0E",x"3E",x"FF",x"32",x"32",x"0E",x"21",x"15",x"0D",x"11",x"26",
x"0D",x"ED",x"53",x"2C",x"0E",x"4E",x"0C",x"06",x"00",x"ED",x"43",x"26",x"0E",x"ED",
x"B0",x"ED",x"53",x"28",x"0E",x"11",x"15",x"0D",x"AF",x"C9",x"EB",x"7E",x"FE",x"11",
x"38",x"02",x"3E",x"10",x"12",x"B7",x"C8",x"47",x"23",x"13",x"7E",x"FE",x"61",x"38",
x"12",x"FE",x"7B",x"30",x"04",x"E6",x"DF",x"18",x"0A",x"FE",x"90",x"38",x"06",x"FE",
x"99",x"30",x"02",x"D6",x"10",x"12",x"10",x"E4",x"C9",x"36",x"00",x"23",x"0B",x"78",
x"B1",x"20",x"F8",x"C9",x"FA",x"85",x"F5",x"CD",x"6B",x"F7",x"28",x"1C",x"21",x"26",
x"0D",x"22",x"2C",x"0E",x"3E",x"FF",x"32",x"2B",x"0E",x"3A",x"2A",x"0E",x"B7",x"20",
x"0B",x"CD",x"72",x"F9",x"38",x"06",x"08",x"CD",x"7C",x"F5",x"08",x"C9",x"AF",x"32",
x"14",x"0D",x"32",x"2A",x"0E",x"18",x"07",x"AF",x"32",x"F3",x"0B",x"32",x"0C",x"0D",
x"21",x"00",x"00",x"22",x"6F",x"0B",x"C9",x"F2",x"53",x"F6",x"CD",x"62",x"F7",x"C8",
x"CD",x"72",x"F7",x"C0",x"ED",x"4B",x"05",x"0D",x"78",x"B1",x"28",x"1B",x"2A",x"07",
x"0D",x"4E",x"23",x"22",x"07",x"0D",x"2A",x"05",x"0D",x"2B",x"22",x"05",x"0D",x"7C",
x"B5",x"20",x"06",x"3A",x"0E",x"0D",x"32",x"6E",x"0B",x"AF",x"C9",x"3A",x"F3",x"0B",
x"3D",x"3E",x"E7",x"C0",x"21",x"00",x"01",x"22",x"09",x"0D",x"21",x"05",x"0C",x"22",
x"10",x"0D",x"22",x"07",x"0D",x"3A",x"0E",x"0D",x"B7",x"3E",x"EC",x"CC",x"7B",x"F7",
x"30",x"0C",x"3A",x"F3",x"0B",x"3D",x"28",x"BE",x"AF",x"37",x"C9",x"32",x"0B",x"0D",
x"21",x"0B",x"0D",x"7E",x"36",x"EC",x"21",x"0E",x"0D",x"36",x"FF",x"21",x"00",x"00",
x"22",x"05",x"0D",x"21",x"6E",x"0B",x"36",x"FF",x"C9",x"CD",x"62",x"F7",x"C8",x"CD",
x"72",x"F7",x"C0",x"3E",x"FF",x"32",x"F1",x"0B",x"3A",x"F3",x"0B",x"3D",x"20",x"27",
x"C5",x"D5",x"CD",x"9E",x"F5",x"69",x"D1",x"C1",x"B7",x"C0",x"1A",x"BD",x"3E",x"E8",
x"C2",x"EB",x"F5",x"13",x"0B",x"78",x"B1",x"20",x"E9",x"C9",x"F2",x"AD",x"F6",x"CD",
x"62",x"F7",x"C8",x"CD",x"72",x"F7",x"C0",x"3A",x"F3",x"0B",x"3D",x"21",x"9E",x"F5",
x"CA",x"6C",x"F2",x"ED",x"53",x"10",x"0D",x"ED",x"43",x"09",x"0D",x"CD",x"D7",x"F5",
x"C3",x"F4",x"F5",x"CD",x"6B",x"F7",x"C8",x"3A",x"2A",x"0E",x"B7",x"3E",x"EC",x"C0",
x"79",x"32",x"2E",x"0E",x"21",x"2F",x"0E",x"7E",x"B7",x"28",x"04",x"35",x"CA",x"89",
x"F6",x"ED",x"5B",x"26",x"0E",x"21",x"00",x"01",x"B7",x"ED",x"52",x"CA",x"89",x"F6",
x"13",x"ED",x"53",x"26",x"0E",x"2A",x"28",x"0E",x"71",x"23",x"22",x"28",x"0E",x"AF",
x"C9",x"21",x"26",x"0D",x"22",x"2C",x"0E",x"CD",x"72",x"F9",x"38",x"05",x"21",x"2A",
x"0E",x"35",x"C9",x"21",x"01",x"00",x"22",x"26",x"0E",x"3A",x"2E",x"0E",x"21",x"26",
x"0D",x"77",x"23",x"22",x"28",x"0E",x"AF",x"37",x"C9",x"CD",x"6B",x"F7",x"C8",x"3A",
x"14",x"0D",x"3D",x"21",x"57",x"F6",x"CA",x"4B",x"F2",x"3A",x"2A",x"0E",x"B7",x"3E",
x"EC",x"C0",x"C5",x"D5",x"21",x"2F",x"0E",x"7E",x"36",x"00",x"B7",x"37",x"C4",x"89",
x"F6",x"D1",x"C1",x"30",x"C1",x"ED",x"43",x"26",x"0E",x"ED",x"53",x"2C",x"0E",x"C3",
x"66",x"F5",x"2E",x"40",x"B7",x"28",x"01",x"29",x"3A",x"6C",x"0B",x"A5",x"28",x"04",
x"3E",x"C0",x"AD",x"6F",x"F3",x"3A",x"12",x"0B",x"B5",x"14",x"15",x"28",x"01",x"AD",
x"D3",x"05",x"32",x"12",x"0B",x"FB",x"C9",x"F3",x"3A",x"12",x"0B",x"E6",x"3F",x"18",
x"F1",x"AF",x"21",x"F0",x"0B",x"11",x"F1",x"0B",x"01",x"44",x"02",x"77",x"ED",x"B0",
x"32",x"6D",x"0B",x"32",x"6E",x"0B",x"21",x"00",x"00",x"22",x"6F",x"0B",x"3E",x"80",
x"32",x"6C",x"0B",x"3A",x"12",x"0B",x"E6",x"3F",x"32",x"12",x"0B",x"D3",x"05",x"C9",
x"46",x"23",x"C5",x"E5",x"4E",x"F7",x"21",x"E1",x"C1",x"10",x"F6",x"C9",x"21",x"41",
x"F7",x"18",x"EF",x"02",x"0D",x"0A",x"09",x"52",x"65",x"61",x"64",x"69",x"6E",x"67",
x"3A",x"20",x"09",x"53",x"65",x"61",x"72",x"63",x"68",x"69",x"6E",x"67",x"09",x"46",
x"6F",x"75",x"6E",x"64",x"3A",x"20",x"20",x"20",x"AF",x"32",x"F1",x"0B",x"3A",x"F3",
x"0B",x"18",x"03",x"3A",x"14",x"0D",x"B7",x"3E",x"E9",x"C9",x"21",x"0B",x"0D",x"7E",
x"B7",x"C8",x"36",x"EC",x"C9",x"ED",x"73",x"33",x"0E",x"AF",x"57",x"CD",x"DE",x"F6",
x"CD",x"7C",x"FA",x"AF",x"32",x"F0",x"0B",x"D9",x"21",x"00",x"00",x"06",x"00",x"D9",
x"3E",x"DC",x"D3",x"04",x"0E",x"00",x"CD",x"3C",x"F9",x"21",x"00",x"00",x"06",x"20",
x"54",x"CD",x"38",x"F9",x"19",x"10",x"FA",x"29",x"29",x"29",x"7C",x"CB",x"15",x"88",
x"57",x"21",x"00",x"04",x"CD",x"38",x"F9",x"D9",x"80",x"47",x"30",x"01",x"23",x"D9",
x"7B",x"92",x"30",x"02",x"ED",x"44",x"FE",x"03",x"30",x"C1",x"2B",x"7C",x"B5",x"20",
x"E7",x"D9",x"29",x"29",x"29",x"29",x"29",x"29",x"7C",x"CB",x"15",x"CE",x"00",x"D9",
x"F5",x"3E",x"88",x"32",x"F0",x"0B",x"3E",x"E8",x"D3",x"04",x"CD",x"3C",x"F9",x"21",
x"00",x"00",x"E5",x"44",x"54",x"E3",x"CD",x"2B",x"F9",x"19",x"19",x"10",x"F8",x"7C",
x"CB",x"15",x"88",x"57",x"E1",x"7C",x"CB",x"15",x"88",x"67",x"6A",x"D1",x"CD",x"2B",
x"F9",x"7D",x"6C",x"67",x"CD",x"2B",x"F9",x"94",x"30",x"07",x"C6",x"02",x"38",x"F3",
x"C3",x"87",x"F7",x"FE",x"04",x"38",x"EC",x"3E",x"DC",x"D3",x"04",x"CD",x"2B",x"F9",
x"FD",x"21",x"00",x"00",x"DD",x"2A",x"10",x"0D",x"CD",x"19",x"F9",x"D9",x"2A",x"6F",
x"0B",x"ED",x"5B",x"09",x"0D",x"D9",x"CD",x"19",x"F9",x"FE",x"6A",x"C2",x"87",x"F7",
x"CD",x"19",x"F9",x"21",x"13",x"0D",x"BE",x"28",x"09",x"7E",x"FE",x"FF",x"CA",x"87",
x"F7",x"C3",x"FD",x"F8",x"32",x"0F",x"0D",x"CD",x"19",x"F9",x"32",x"F3",x"0B",x"CD",
x"19",x"F9",x"32",x"0C",x"0D",x"CD",x"19",x"F9",x"47",x"C5",x"18",x"06",x"C5",x"D9",
x"2A",x"6F",x"0B",x"D9",x"CD",x"19",x"F9",x"21",x"0D",x"0D",x"BE",x"C2",x"FD",x"F8",
x"CD",x"19",x"F9",x"47",x"CD",x"19",x"F9",x"08",x"D9",x"7A",x"B3",x"1B",x"D9",x"CA",
x"01",x"F9",x"3A",x"F3",x"0B",x"3D",x"28",x"0F",x"3A",x"F1",x"0B",x"B7",x"28",x"09",
x"08",x"DD",x"BE",x"00",x"28",x"07",x"C3",x"09",x"F9",x"08",x"DD",x"77",x"00",x"DD",
x"23",x"FD",x"23",x"10",x"D5",x"CD",x"19",x"F9",x"32",x"0E",x"0D",x"D9",x"E5",x"D9",
x"CD",x"19",x"F9",x"BF",x"08",x"E1",x"44",x"CD",x"19",x"F9",x"4D",x"67",x"08",x"6F",
x"ED",x"42",x"C1",x"20",x"40",x"FD",x"22",x"05",x"0D",x"DD",x"22",x"10",x"0D",x"21",
x"0D",x"0D",x"34",x"D9",x"ED",x"53",x"09",x"0D",x"D9",x"10",x"91",x"3A",x"F3",x"0B",
x"3D",x"28",x"0C",x"3A",x"13",x"0D",x"FE",x"FF",x"28",x"05",x"D9",x"7A",x"B3",x"20",
x"1E",x"C3",x"BD",x"FA",x"3E",x"F5",x"32",x"2A",x"0E",x"18",x"05",x"3E",x"F5",x"32",
x"0B",x"0D",x"21",x"62",x"0B",x"CB",x"DE",x"06",x"00",x"10",x"FE",x"18",x"11",x"3E",
x"EA",x"18",x"0A",x"3A",x"F1",x"0B",x"B7",x"3E",x"E7",x"28",x"02",x"3E",x"E8",x"32",
x"0B",x"0D",x"F5",x"CD",x"BD",x"FA",x"F1",x"B7",x"ED",x"7B",x"33",x"0E",x"C9",x"26",
x"80",x"CD",x"38",x"F9",x"BA",x"F5",x"9F",x"CD",x"F7",x"FA",x"F1",x"CB",x"1C",x"30",
x"F2",x"7C",x"C9",x"DB",x"59",x"E6",x"20",x"EE",x"20",x"4F",x"1E",x"00",x"FB",x"76",
x"18",x"0F",x"1E",x"00",x"FB",x"76",x"1C",x"CC",x"69",x"F9",x"DB",x"59",x"A9",x"E6",
x"20",x"28",x"F5",x"1C",x"CC",x"69",x"F9",x"DB",x"59",x"A9",x"E6",x"20",x"20",x"F5",
x"DB",x"5B",x"D3",x"07",x"3A",x"F0",x"0B",x"B7",x"28",x"0D",x"FE",x"88",x"3E",x"A0",
x"28",x"02",x"3E",x"88",x"32",x"F0",x"0B",x"D3",x"00",x"DB",x"58",x"E6",x"18",x"CA",
x"ED",x"F8",x"7B",x"C9",x"ED",x"73",x"33",x"0E",x"AF",x"57",x"3D",x"CD",x"DE",x"F6",
x"01",x"00",x"00",x"E3",x"0B",x"78",x"B1",x"20",x"FA",x"CD",x"7C",x"FA",x"3E",x"88",
x"32",x"F0",x"0B",x"01",x"14",x"00",x"3A",x"32",x"0E",x"B7",x"28",x"03",x"01",x"28",
x"00",x"CD",x"31",x"FA",x"CD",x"62",x"FA",x"CD",x"62",x"FA",x"CD",x"3D",x"FA",x"2A",
x"6F",x"0B",x"D9",x"0E",x"6A",x"CD",x"3D",x"FA",x"FD",x"2A",x"2C",x"0E",x"3A",x"32",
x"0E",x"4F",x"CD",x"3D",x"FA",x"3A",x"14",x"0D",x"4F",x"CD",x"3D",x"FA",x"3A",x"30",
x"0E",x"4F",x"CD",x"3D",x"FA",x"2A",x"26",x"0E",x"4C",x"7D",x"B7",x"28",x"01",x"0C",
x"CD",x"3D",x"FA",x"18",x"05",x"D9",x"2A",x"6F",x"0B",x"D9",x"3A",x"31",x"0E",x"4F",
x"CD",x"3D",x"FA",x"7C",x"B7",x"55",x"28",x"02",x"AF",x"57",x"4A",x"CD",x"3D",x"FA",
x"FD",x"4E",x"00",x"FD",x"23",x"2B",x"CD",x"3D",x"FA",x"15",x"20",x"F4",x"7C",x"B5",
x"3A",x"2B",x"0E",x"28",x"01",x"AF",x"4F",x"CD",x"3D",x"FA",x"EB",x"D9",x"4D",x"CD",
x"3D",x"FA",x"4C",x"CD",x"3D",x"FA",x"D9",x"EB",x"22",x"26",x"0E",x"FD",x"22",x"2C",
x"0E",x"3A",x"31",x"0E",x"3C",x"32",x"31",x"0E",x"7C",x"B5",x"20",x"B3",x"01",x"01",
x"05",x"CD",x"31",x"FA",x"FB",x"76",x"AF",x"32",x"32",x"0E",x"C3",x"BD",x"FA",x"CD",
x"5D",x"FA",x"CD",x"5D",x"FA",x"10",x"F8",x"0D",x"20",x"F5",x"C9",x"06",x"08",x"CB",
x"09",x"CD",x"4F",x"FA",x"CB",x"79",x"CD",x"F7",x"FA",x"CD",x"4F",x"FA",x"10",x"F1",
x"C9",x"CB",x"79",x"28",x"05",x"3A",x"F4",x"FA",x"18",x"0D",x"3A",x"F5",x"FA",x"18",
x"08",x"3A",x"F3",x"FA",x"18",x"03",x"3A",x"F6",x"FA",x"08",x"DB",x"58",x"E6",x"18",
x"CA",x"E6",x"F8",x"FB",x"76",x"D3",x"50",x"08",x"D3",x"04",x"DB",x"5B",x"D3",x"07",
x"CD",x"56",x"F9",x"C9",x"F3",x"AF",x"D3",x"58",x"D3",x"59",x"D3",x"5A",x"D3",x"5B",
x"D3",x"04",x"3D",x"32",x"71",x"0B",x"3A",x"11",x"0B",x"E6",x"F0",x"F6",x"07",x"D3",
x"03",x"3A",x"12",x"0B",x"E6",x"EF",x"32",x"12",x"0B",x"E6",x"C0",x"F6",x"2F",x"D3",
x"05",x"AF",x"32",x"14",x"0B",x"3E",x"0A",x"D3",x"70",x"3E",x"23",x"D3",x"71",x"DB",
x"5B",x"D3",x"07",x"21",x"38",x"00",x"7E",x"36",x"C9",x"32",x"F2",x"0B",x"C9",x"F3",
x"CD",x"FF",x"F6",x"3A",x"11",x"0B",x"D3",x"03",x"3A",x"12",x"0B",x"D3",x"05",x"3A",
x"1F",x"0B",x"47",x"CB",x"40",x"28",x"08",x"3E",x"0A",x"D3",x"70",x"3E",x"03",x"D3",
x"71",x"78",x"07",x"07",x"D3",x"5B",x"07",x"D3",x"5A",x"07",x"D3",x"59",x"07",x"D3",
x"58",x"3A",x"F2",x"0B",x"32",x"38",x"00",x"AF",x"37",x"FB",x"C9",x"D6",x"DE",x"CE",
x"BC",x"D9",x"3E",x"80",x"20",x"01",x"AF",x"AC",x"17",x"30",x"09",x"7C",x"EE",x"08",
x"67",x"7D",x"EE",x"10",x"6F",x"37",x"ED",x"6A",x"D9",x"C9",x"FF",x"01",x"02",x"FF",
x"FF",x"05",x"06",x"FF",x"00",x"FF",x"02",x"FF",x"04",x"05",x"06",x"FF",x"C3",x"23",
x"0B",x"00",x"00",x"00",x"00",x"00",x"F5",x"3E",x"70",x"D3",x"02",x"C3",x"12",x"C4",
x"E3",x"7E",x"23",x"E3",x"08",x"F5",x"3A",x"03",x"00",x"F5",x"3E",x"70",x"32",x"03",
x"00",x"D3",x"02",x"C3",x"63",x"C3",x"08",x"F1",x"32",x"03",x"00",x"D3",x"02",x"F1",
x"08",x"C9",x"32",x"03",x"00",x"D3",x"02",x"F1",x"FB",x"C9",x"4D",x"4F",x"50",x"53",
x"03",x"56",x"47",x"42",x"05",x"52",x"53",x"32",x"33",x"32",x"04",x"44",x"49",x"53",
x"4B",x"43",x"49",x"53",x"4C",x"08",x"08",x"3E",x"6B",x"63",x"7F",x"63",x"63",x"00",
x"00",x"08",x"08",x"7E",x"68",x"60",x"7C",x"60",x"7E",x"00",x"00",x"08",x"08",x"3C",
x"18",x"18",x"18",x"18",x"3C",x"00",x"00",x"08",x"08",x"3E",x"6B",x"63",x"63",x"63",
x"3E",x"00",x"00",x"14",x"00",x"3E",x"63",x"63",x"63",x"63",x"3E",x"00",x"00",x"14",
x"14",x"3E",x"63",x"63",x"63",x"63",x"3E",x"00",x"00",x"08",x"08",x"6B",x"63",x"63",
x"63",x"63",x"3E",x"00",x"00",x"14",x"00",x"63",x"63",x"63",x"63",x"63",x"3E",x"00",
x"00",x"14",x"14",x"77",x"63",x"63",x"63",x"63",x"3E",x"00",x"00",x"00",x"00",x"00",
x"00",x"1F",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1F",x"1F",x"00",
x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"1F",x"1F",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"00",x"FF",
x"FF",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",
x"18",x"FF",x"E7",x"C3",x"99",x"99",x"81",x"99",x"99",x"FF",x"FF",x"08",x"08",x"08",
x"3C",x"06",x"3E",x"66",x"3E",x"00",x"00",x"08",x"08",x"08",x"3C",x"66",x"7E",x"60",
x"3C",x"00",x"00",x"08",x"08",x"00",x"38",x"18",x"18",x"18",x"3C",x"00",x"00",x"08",
x"08",x"08",x"3C",x"66",x"66",x"66",x"3C",x"00",x"00",x"00",x"24",x"00",x"3C",x"66",
x"66",x"66",x"3C",x"00",x"00",x"24",x"24",x"00",x"3C",x"66",x"66",x"66",x"3C",x"00",
x"00",x"08",x"08",x"08",x"66",x"66",x"66",x"66",x"3E",x"00",x"00",x"00",x"24",x"00",
x"66",x"66",x"66",x"66",x"3E",x"00",x"00",x"24",x"24",x"00",x"66",x"66",x"66",x"66",
x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"F8",x"F8",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"18",x"F8",x"F8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
x"FF",x"00",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"F8",x"F8",x"18",x"18",x"18",
x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"C3",x"99",
x"9F",x"9F",x"9F",x"99",x"C3",x"FF",x"FF",x"FF",x"C3",x"99",x"9F",x"C3",x"F9",x"99",
x"C3",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D9",
x"C5",x"D5",x"E5",x"2A",x"2E",x"17",x"E5",x"FD",x"E3",x"AF",x"47",x"4F",x"D9",x"67",
x"6F",x"57",x"5F",x"47",x"4F",x"FD",x"7E",x"00",x"FD",x"23",x"E5",x"C5",x"21",x"3F",
x"FF",x"01",x"0B",x"00",x"ED",x"B1",x"20",x"6B",x"CB",x"21",x"21",x"4A",x"FF",x"09",
x"7E",x"23",x"66",x"6F",x"C1",x"E3",x"7D",x"B7",x"C9",x"3E",x"40",x"DA",x"3E",x"80",
x"20",x"57",x"F5",x"B1",x"4F",x"F1",x"EE",x"03",x"A1",x"4F",x"18",x"CF",x"20",x"4B",
x"CB",x"C9",x"18",x"C9",x"20",x"45",x"2C",x"18",x"C4",x"2C",x"24",x"D9",x"78",x"B1",
x"D9",x"20",x"BC",x"25",x"FD",x"7E",x"FF",x"FE",x"2A",x"5F",x"28",x"B3",x"1E",x"30",
x"18",x"AF",x"3E",x"04",x"21",x"5C",x"FD",x"C3",x"F0",x"FF",x"2C",x"D9",x"78",x"B1",
x"D9",x"28",x"A0",x"24",x"18",x"9D",x"D9",x"78",x"B1",x"20",x"04",x"FD",x"E5",x"C1",
x"0B",x"D9",x"14",x"18",x"90",x"D9",x"78",x"B1",x"20",x"DC",x"FD",x"E5",x"C1",x"0B",
x"D9",x"18",x"84",x"C1",x"E1",x"D9",x"78",x"B1",x"20",x"04",x"FD",x"E5",x"C1",x"0B",
x"FD",x"E1",x"D9",x"22",x"1C",x"17",x"7A",x"FE",x"04",x"30",x"0D",x"B7",x"C2",x"1A",
x"FD",x"FD",x"7E",x"08",x"E6",x"7F",x"D6",x"3F",x"84",x"6F",x"C5",x"FD",x"7E",x"06",
x"B7",x"28",x"11",x"FD",x"7E",x"08",x"E6",x"80",x"28",x"0A",x"FD",x"AE",x"08",x"FD",
x"77",x"08",x"C1",x"CB",x"C1",x"3E",x"C1",x"FD",x"7E",x"08",x"D6",x"3F",x"47",x"D9",
x"59",x"50",x"D9",x"AF",x"67",x"6F",x"B2",x"20",x"05",x"B0",x"FA",x"96",x"FD",x"68",
x"D9",x"1B",x"B7",x"ED",x"52",x"19",x"1A",x"D9",x"28",x"02",x"30",x"19",x"FE",x"2C",
x"28",x"01",x"37",x"14",x"15",x"20",x"0B",x"2C",x"2D",x"FA",x"B8",x"FD",x"28",x"06",
x"30",x"E2",x"2D",x"B7",x"30",x"DE",x"24",x"18",x"DB",x"CB",x"49",x"28",x"01",x"25",
x"CB",x"41",x"20",x"05",x"79",x"E6",x"FC",x"28",x"01",x"25",x"CB",x"7C",x"C2",x"1A",
x"FD",x"7D",x"3D",x"F2",x"1A",x"FD",x"14",x"15",x"20",x"14",x"AF",x"CB",x"78",x"20",
x"01",x"78",x"6F",x"B7",x"20",x"0E",x"24",x"25",x"28",x"0A",x"CB",x"D1",x"2E",x"01",
x"18",x"04",x"6C",x"78",x"94",x"47",x"14",x"15",x"20",x"06",x"1C",x"1D",x"20",x"02",
x"1E",x"20",x"C4",x"62",x"FF",x"24",x"25",x"28",x"13",x"14",x"15",x"20",x"0F",x"CB",
x"51",x"28",x"05",x"7C",x"3D",x"CC",x"60",x"FF",x"7B",x"CD",x"8D",x"FF",x"18",x"EA",
x"7B",x"FE",x"20",x"CC",x"62",x"FF",x"D9",x"59",x"50",x"D9",x"04",x"05",x"28",x"03",
x"F2",x"29",x"FE",x"7D",x"3D",x"28",x"16",x"2C",x"2D",x"28",x"12",x"D9",x"1B",x"1A",
x"FE",x"2C",x"28",x"FA",x"D9",x"18",x"F3",x"CD",x"96",x"FF",x"06",x"04",x"48",x"18",
x"33",x"D5",x"48",x"C5",x"58",x"1D",x"FD",x"7E",x"08",x"D6",x"3B",x"4F",x"D6",x"04",
x"2A",x"1C",x"17",x"25",x"84",x"FA",x"37",x"FE",x"BC",x"30",x"03",x"7C",x"0E",x"04",
x"C6",x"04",x"47",x"68",x"05",x"78",x"FE",x"10",x"3E",x"00",x"DC",x"87",x"FF",x"B7",
x"20",x"08",x"78",x"3D",x"B9",x"30",x"EF",x"2E",x"00",x"D2",x"48",x"0C",x"06",x"04",
x"D9",x"EB",x"B7",x"ED",x"42",x"09",x"EB",x"28",x"17",x"1A",x"13",x"D9",x"FE",x"2C",
x"28",x"0B",x"78",x"FE",x"10",x"3E",x"00",x"DC",x"87",x"FF",x"C6",x"30",x"04",x"CD",
x"8D",x"FF",x"18",x"E0",x"0A",x"FE",x"2E",x"20",x"45",x"CD",x"8D",x"FF",x"03",x"0A",
x"FE",x"2C",x"28",x"F7",x"D9",x"7A",x"B7",x"20",x"0C",x"3A",x"1D",x"17",x"2F",x"BB",
x"30",x"05",x"AF",x"1C",x"FA",x"DB",x"FE",x"D9",x"0A",x"FE",x"2A",x"28",x"0B",x"FE",
x"25",x"28",x"07",x"FE",x"23",x"20",x"1D",x"D9",x"18",x"0C",x"D9",x"78",x"91",x"38",
x"07",x"B5",x"28",x"0C",x"3E",x"F0",x"18",x"08",x"78",x"FE",x"10",x"3E",x"00",x"DC",
x"87",x"FF",x"04",x"D9",x"C6",x"30",x"18",x"BB",x"0A",x"FE",x"5E",x"D9",x"C1",x"D1",
x"41",x"20",x"47",x"FD",x"7E",x"06",x"B7",x"20",x"01",x"47",x"3E",x"45",x"CD",x"8D",
x"FF",x"CB",x"78",x"3E",x"2B",x"28",x"06",x"78",x"ED",x"44",x"47",x"3E",x"2D",x"CD",
x"8D",x"FF",x"15",x"7A",x"FE",x"04",x"38",x"0A",x"3E",x"30",x"CD",x"8D",x"FF",x"D9",
x"03",x"D9",x"18",x"F0",x"78",x"01",x"FF",x"0A",x"90",x"0C",x"30",x"FC",x"80",x"47",
x"79",x"C6",x"30",x"CD",x"8D",x"FF",x"78",x"C6",x"30",x"CD",x"8D",x"FF",x"D9",x"03",
x"03",x"03",x"03",x"D9",x"D9",x"ED",x"43",x"2E",x"17",x"E1",x"D1",x"C1",x"D9",x"21",
x"7A",x"E6",x"C3",x"F0",x"FF",x"2B",x"2D",x"24",x"3C",x"3E",x"2A",x"25",x"23",x"2C",
x"5E",x"2E",x"39",x"FD",x"2C",x"FD",x"C9",x"FC",x"22",x"FD",x"05",x"FD",x"05",x"FD",
x"00",x"FD",x"00",x"FD",x"FA",x"FC",x"EC",x"FC",x"E9",x"FC",x"1E",x"30",x"CB",x"49",
x"3E",x"24",x"C4",x"8D",x"FF",x"CB",x"41",x"3E",x"2D",x"20",x"1E",x"79",x"E6",x"F8",
x"87",x"3E",x"20",x"38",x"16",x"F0",x"3E",x"2B",x"18",x"11",x"3D",x"F8",x"F5",x"3E",
x"20",x"CD",x"8D",x"FF",x"F1",x"18",x"F5",x"E5",x"21",x"CE",x"F7",x"18",x"04",x"E5",
x"21",x"B3",x"FE",x"CD",x"F0",x"FF",x"E1",x"C9",x"21",x"14",x"FA",x"C3",x"F0",x"FF",
x"2A",x"2E",x"17",x"7E",x"11",x"00",x"00",x"FE",x"3C",x"28",x"06",x"1C",x"FE",x"3E",
x"20",x"06",x"1C",x"14",x"23",x"22",x"2E",x"17",x"7E",x"FE",x"23",x"28",x"F6",x"FE",
x"25",x"28",x"F2",x"FE",x"2A",x"28",x"EE",x"FD",x"7E",x"01",x"92",x"ED",x"44",x"FA",
x"1A",x"FD",x"1D",x"FA",x"D2",x"FF",x"4F",x"20",x"02",x"CB",x"39",x"91",x"F5",x"79",
x"F4",x"7C",x"FF",x"F1",x"21",x"4F",x"E6",x"C3",x"F0",x"FF",x"28",x"43",x"29",x"31",
x"39",x"38",x"35",x"49",x"53",x"4C",x"3E",x"04",x"C3",x"9C",x"F2",x"00",x"00",x"00",
x"F5",x"3E",x"70",x"32",x"03",x"00",x"D3",x"02",x"F1",x"E9",x"7B",x"E6",x"1F",x"1B",
x"FE",x"04"
  );

signal  do : std_logic_vector(7 downto 0);

begin

  process(CLK)
  begin
    if rising_edge(CLK) then
	   do <= myROM(conv_integer(A));
	 end if;
  end process;  
  DOUT <= do;
  
end Behavioral;
