----------------------------------------------------------------------------------
-- Engineer: Jozsef Laszlo ( rbendr AT gmail DOT com )
-- 
-- Create Date:    08:47:30 03/05/2017 
-- Design Name: 	 TVC main rom
-- Module Name:    soundctrl - Behavioral 
-- Project Name:   TVC Home computer VHDL version
-- Description: 
--		rom dumped from TVC emulator
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: All rights reserved
-- Status: works
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity rom16k is
    Port ( CLK : in  STD_LOGIC;
             A : in  STD_LOGIC_VECTOR (13 downto 0);
          DOUT : out STD_LOGIC_VECTOR (7 downto 0)
		   );
				
end rom16k;

architecture Behavioral of rom16k is

type  
  romarray is array(0 to 16383) of std_logic_vector(7 downto 0);

constant
  myROM : romarray := (

--x"F3",x"31",x"FF",x"7F",x"C3",x"80",x"00",x"00",x"ED",x"4D",x"00",x"00",x"00",x"00",
--x"00",x"00",x"ED",x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"ED",x"4D",x"00",x"00",
--x"00",x"00",x"00",x"00",x"ED",x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"ED",x"4D",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--x"E5",x"2A",x"02",x"40",x"E5",x"C9",x"E1",x"ED",x"4D",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"00",x"00",x"E5",x"2A",x"00",x"40",x"E5",x"C9",x"E1",x"ED",x"45",x"00",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"CD",x"7B",x"03",x"C3",x"E0",x"03",x"00",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--x"00",x"00",x"00",x"00",x"00",x"00",x"C5",x"D5",x"E5",x"21",x"00",x"80",x"11",x"01",
--x"80",x"01",x"FF",x"3B",x"75",x"ED",x"B0",x"E1",x"D1",x"C1",x"C9",x"01",x"D7",x"00",
--x"1E",x"00",x"7B",x"D3",x"70",x"6B",x"26",x"00",x"09",x"7E",x"D3",x"71",x"1C",x"7B",
--x"D6",x"10",x"38",x"F0",x"C9",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"77",
--x"BB",x"DD",x"EE",x"55",x"AA",x"63",x"40",x"4B",x"32",x"4D",x"02",x"3C",x"42",x"00",
--x"03",x"03",x"03",x"00",x"00",x"0E",x"FF",x"DD",x"E5",x"DD",x"21",x"00",x"00",x"DD",
--x"39",x"DD",x"7E",x"04",x"E6",x"07",x"5F",x"DD",x"6E",x"06",x"DD",x"66",x"07",x"29",
--x"29",x"29",x"29",x"29",x"29",x"01",x"00",x"80",x"09",x"DD",x"4E",x"04",x"DD",x"46",
--x"05",x"CB",x"38",x"CB",x"19",x"CB",x"38",x"CB",x"19",x"CB",x"38",x"CB",x"19",x"09",
--x"4D",x"44",x"0A",x"57",x"7B",x"C6",x"C9",x"6F",x"3E",x"00",x"CE",x"00",x"67",x"7E",
--x"B2",x"02",x"DD",x"E1",x"C9",x"DD",x"E5",x"DD",x"21",x"00",x"00",x"DD",x"39",x"DD",
--x"7E",x"04",x"E6",x"03",x"5F",x"DD",x"6E",x"06",x"DD",x"66",x"07",x"29",x"29",x"29",
--x"29",x"29",x"29",x"01",x"00",x"80",x"09",x"DD",x"4E",x"04",x"DD",x"46",x"05",x"CB",
--x"38",x"CB",x"19",x"CB",x"38",x"CB",x"19",x"09",x"4D",x"44",x"0A",x"57",x"3E",x"D1",
--x"83",x"6F",x"3E",x"00",x"CE",x"00",x"67",x"7E",x"A2",x"57",x"2E",x"00",x"DD",x"CB",
--x"08",x"46",x"28",x"02",x"2E",x"08",x"DD",x"CB",x"08",x"4E",x"28",x"02",x"CB",x"FD",
--x"1C",x"18",x"02",x"CB",x"3D",x"1D",x"20",x"FB",x"7A",x"B5",x"02",x"DD",x"E1",x"C9",
--x"DD",x"E5",x"DD",x"21",x"00",x"00",x"DD",x"39",x"DD",x"7E",x"04",x"E6",x"01",x"5F",
--x"DD",x"6E",x"06",x"DD",x"66",x"07",x"29",x"29",x"29",x"29",x"29",x"29",x"01",x"00",
--x"80",x"09",x"DD",x"4E",x"04",x"DD",x"46",x"05",x"CB",x"38",x"CB",x"19",x"09",x"4D",
--x"44",x"0A",x"57",x"3E",x"D5",x"83",x"6F",x"3E",x"00",x"CE",x"00",x"67",x"7E",x"A2",
--x"57",x"2E",x"00",x"DD",x"CB",x"08",x"46",x"28",x"02",x"2E",x"02",x"DD",x"CB",x"08",
--x"4E",x"28",x"02",x"CB",x"DD",x"DD",x"CB",x"08",x"56",x"28",x"02",x"CB",x"ED",x"DD",
--x"CB",x"08",x"5E",x"28",x"02",x"CB",x"FD",x"1C",x"18",x"02",x"CB",x"3D",x"1D",x"20",
--x"FB",x"7A",x"B5",x"02",x"DD",x"E1",x"C9",x"3E",x"00",x"D3",x"06",x"CD",x"A0",x"00",
--x"01",x"00",x"00",x"C5",x"21",x"00",x"00",x"E5",x"C5",x"CD",x"E7",x"00",x"F1",x"F1",
--x"C1",x"C5",x"21",x"EF",x"00",x"E5",x"C5",x"CD",x"E7",x"00",x"F1",x"F1",x"C1",x"03",
--x"78",x"D6",x"02",x"38",x"E2",x"01",x"00",x"00",x"C5",x"C5",x"21",x"00",x"00",x"E5",
--x"CD",x"E7",x"00",x"F1",x"F1",x"C1",x"C5",x"C5",x"21",x"FF",x"01",x"E5",x"CD",x"E7",
--x"00",x"F1",x"F1",x"C1",x"03",x"79",x"D6",x"F0",x"78",x"DE",x"00",x"38",x"DF",x"01",
--x"00",x"00",x"C5",x"C5",x"C5",x"CD",x"E7",x"00",x"F1",x"F1",x"C1",x"3E",x"FF",x"91",
--x"5F",x"3E",x"01",x"98",x"57",x"C5",x"D5",x"C5",x"D5",x"CD",x"E7",x"00",x"F1",x"F1",
--x"D1",x"C1",x"3E",x"EF",x"91",x"6F",x"3E",x"00",x"98",x"67",x"E5",x"C5",x"D5",x"E5",
--x"C5",x"CD",x"E7",x"00",x"F1",x"F1",x"D1",x"C1",x"E1",x"C5",x"E5",x"D5",x"CD",x"E7",
--x"00",x"F1",x"F1",x"C1",x"03",x"79",x"D6",x"F0",x"78",x"DE",x"00",x"38",x"BD",x"C9",
--x"3E",x"01",x"D3",x"06",x"CD",x"A0",x"00",x"01",x"00",x"00",x"C5",x"3E",x"01",x"F5",
--x"33",x"21",x"00",x"00",x"E5",x"C5",x"CD",x"2B",x"01",x"F1",x"F1",x"33",x"C1",x"C5",
--x"3E",x"01",x"F5",x"33",x"21",x"EF",x"00",x"E5",x"C5",x"CD",x"2B",x"01",x"F1",x"F1",
--x"33",x"C1",x"03",x"78",x"D6",x"01",x"38",x"D8",x"01",x"00",x"00",x"C5",x"3E",x"02",
--x"F5",x"33",x"C5",x"21",x"00",x"00",x"E5",x"CD",x"2B",x"01",x"F1",x"F1",x"33",x"C1",
--x"C5",x"3E",x"03",x"F5",x"33",x"C5",x"21",x"FF",x"00",x"E5",x"CD",x"2B",x"01",x"F1",
--x"F1",x"33",x"C1",x"03",x"79",x"D6",x"F0",x"78",x"DE",x"00",x"38",x"D5",x"01",x"00",
--x"00",x"51",x"C5",x"D5",x"33",x"C5",x"C5",x"CD",x"2B",x"01",x"F1",x"F1",x"33",x"C1",
--x"03",x"79",x"D6",x"F0",x"78",x"DE",x"00",x"38",x"EA",x"C9",x"3E",x"02",x"D3",x"06",
--x"CD",x"A0",x"00",x"01",x"00",x"00",x"C5",x"3E",x"0F",x"F5",x"33",x"21",x"00",x"00",
--x"E5",x"C5",x"CD",x"88",x"01",x"F1",x"F1",x"33",x"C1",x"C5",x"3E",x"0F",x"F5",x"33",
--x"21",x"EF",x"00",x"E5",x"C5",x"CD",x"88",x"01",x"F1",x"F1",x"33",x"C1",x"03",x"79",
--x"D6",x"7F",x"78",x"DE",x"00",x"38",x"D5",x"01",x"00",x"00",x"C5",x"3E",x"0F",x"F5",
--x"33",x"C5",x"21",x"00",x"00",x"E5",x"CD",x"88",x"01",x"F1",x"F1",x"33",x"C1",x"C5",
--x"3E",x"0F",x"F5",x"33",x"C5",x"21",x"7F",x"00",x"E5",x"CD",x"88",x"01",x"F1",x"F1",
--x"33",x"C1",x"03",x"79",x"D6",x"F0",x"78",x"DE",x"00",x"38",x"D5",x"01",x"00",x"00",
--x"51",x"C5",x"D5",x"33",x"C5",x"C5",x"CD",x"88",x"01",x"F1",x"F1",x"33",x"C1",x"03",
--x"79",x"D6",x"7F",x"78",x"DE",x"00",x"38",x"EA",x"C9",x"DD",x"E5",x"DD",x"21",x"00",
--x"00",x"DD",x"39",x"F5",x"3E",x"00",x"D3",x"06",x"CD",x"B3",x"00",x"0E",x"00",x"11",
--x"00",x"00",x"79",x"B7",x"20",x"07",x"C5",x"D5",x"CD",x"F1",x"01",x"D1",x"C1",x"79",
--x"3D",x"20",x"07",x"C5",x"D5",x"CD",x"84",x"02",x"D1",x"C1",x"79",x"D6",x"02",x"20",
--x"07",x"C5",x"D5",x"CD",x"FE",x"02",x"D1",x"C1",x"0C",x"79",x"D6",x"03",x"20",x"01",
--x"4F",x"06",x"00",x"7B",x"E6",x"01",x"D3",x"A0",x"13",x"21",x"10",x"27",x"E3",x"00",
--x"DD",x"6E",x"FE",x"DD",x"66",x"FF",x"2B",x"33",x"33",x"E5",x"7C",x"B5",x"20",x"F1",
--x"04",x"78",x"D6",x"20",x"38",x"E1",x"18",x"B4",x"3E",x"02",x"CF",x"C9",x"3E",x"00",
--x"CF",x"76",x"18",x"FD",
--      
--x"f3",x"31",x"ff",x"7f",x"21",x"3c",x"00",x"06",x"10",x"0e",x"00",x"79",x"d3",x"70",x"7e",x"d3",
--x"71",x"0c",x"23",x"10",x"f6",x"dd",x"21",x"3f",x"80",x"21",x"00",x"80",x"11",x"40",x"00",x"06",
--x"f0",x"3e",x"80",x"77",x"dd",x"36",x"00",x"01",x"19",x"dd",x"19",x"10",x"f6",x"7b",x"d3",x"a0",
--x"1c",x"01",x"30",x"75",x"00",x"0b",x"78",x"b1",x"20",x"fa",x"18",x"f1",x"63",x"40",x"4b",x"32",
--x"4d",x"02",x"3c",x"42",x"00",x"03",x"03",x"03",x"00",x"00",x"0e",x"ff",x"00",x"00",x"00",x"00",
--
--x"f3",x"31",x"ff",x"7f",x"21",x"24",x"00",x"06",x"10",x"0e",x"00",x"79",x"d3",x"70",x"7e",x"d3",
--x"71",x"0c",x"23",x"10",x"f6",x"7b",x"d3",x"a0",x"1c",x"01",x"30",x"75",x"00",x"0b",x"78",x"b1",
--x"20",x"fa",x"18",x"f1",x"63",x"40",x"4c",x"32",x"4d",x"02",x"3c",x"42",x"00",x"03",x"03",x"03",
--x"00",x"00",x"0e",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

--others => x"ff"


-- TVC ORIGINAL ROM DUMP
x"C3",x"29",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"01",x"02",x"03",x"04",x"05",x"06",x"07",x"08",x"09",x"00",x"02",x"04",x"06",x"08",
x"10",x"12",x"14",x"16",x"18",x"00",x"03",x"06",x"09",x"12",x"15",x"18",x"21",x"24",
x"27",x"00",x"04",x"08",x"12",x"16",x"20",x"24",x"28",x"32",x"36",x"00",x"05",x"10",
x"15",x"20",x"25",x"30",x"35",x"40",x"45",x"00",x"06",x"12",x"18",x"24",x"30",x"36",
x"42",x"48",x"54",x"00",x"07",x"14",x"21",x"28",x"35",x"42",x"49",x"56",x"63",x"00",
x"08",x"16",x"24",x"32",x"40",x"48",x"56",x"64",x"72",x"00",x"09",x"18",x"27",x"36",
x"45",x"54",x"63",x"72",x"81",x"BB",x"DB",x"BB",x"DB",x"80",x"DB",x"BB",x"DB",x"F2",
x"DF",x"9B",x"E8",x"FC",x"DF",x"65",x"DD",x"02",x"E0",x"93",x"DD",x"53",x"E0",x"04",
x"E1",x"0E",x"E1",x"5C",x"E1",x"10",x"E9",x"82",x"E3",x"B2",x"E3",x"33",x"E7",x"EE",
x"E2",x"CB",x"E1",x"C1",x"E3",x"85",x"DD",x"80",x"DD",x"51",x"E9",x"52",x"E4",x"08",
x"DE",x"B6",x"E4",x"06",x"DB",x"32",x"E3",x"C9",x"E8",x"73",x"E5",x"42",x"E5",x"54",
x"E7",x"53",x"E5",x"73",x"E5",x"C7",x"E6",x"1B",x"E2",x"F4",x"E6",x"0F",x"E7",x"1B",
x"DE",x"82",x"E9",x"90",x"E7",x"33",x"E8",x"A3",x"FF",x"31",x"DE",x"D3",x"E9",x"17",
x"E1",x"70",x"E5",x"93",x"F4",x"FB",x"F5",x"12",x"F5",x"8E",x"F4",x"26",x"F7",x"82",
x"EA",x"9F",x"EA",x"9A",x"EA",x"D2",x"EA",x"CD",x"EA",x"C3",x"EA",x"BE",x"EA",x"92",
x"FA",x"28",x"FB",x"68",x"EA",x"43",x"6F",x"70",x"79",x"72",x"69",x"67",x"68",x"74",
x"20",x"28",x"63",x"29",x"20",x"31",x"39",x"38",x"34",x"20",x"20",x"49",x"6E",x"74",
x"65",x"6C",x"6C",x"69",x"67",x"65",x"6E",x"74",x"20",x"53",x"6F",x"66",x"74",x"77",
x"61",x"72",x"65",x"20",x"4C",x"74",x"64",x"00",x"00",x"00",x"00",x"00",x"50",x"3F",
x"00",x"00",x"00",x"00",x"00",x"10",x"40",x"31",x"24",x"19",x"49",x"79",x"26",x"3F",
x"57",x"07",x"08",x"05",x"32",x"17",x"40",x"69",x"75",x"80",x"50",x"20",x"73",x"3F",
x"74",x"48",x"34",x"08",x"40",x"14",x"C0",x"98",x"88",x"84",x"26",x"00",x"72",x"BF",
x"19",x"89",x"03",x"25",x"20",x"43",x"40",x"99",x"45",x"58",x"22",x"52",x"47",x"40",
x"07",x"38",x"96",x"88",x"85",x"86",x"3F",x"00",x"00",x"00",x"00",x"51",x"11",x"40",
x"23",x"70",x"49",x"46",x"25",x"29",x"3C",x"06",x"95",x"88",x"64",x"44",x"50",x"42",
x"63",x"75",x"99",x"82",x"00",x"14",x"41",x"16",x"65",x"64",x"73",x"28",x"33",x"3E",
x"01",x"79",x"97",x"92",x"08",x"10",x"43",x"97",x"10",x"08",x"94",x"20",x"11",x"42",
x"99",x"92",x"50",x"58",x"02",x"23",x"40",x"90",x"37",x"14",x"68",x"15",x"29",x"C0",
x"57",x"15",x"49",x"03",x"63",x"31",x"40",x"78",x"14",x"60",x"81",x"35",x"67",x"BF",
x"42",x"95",x"06",x"04",x"07",x"10",x"C1",x"21",x"40",x"81",x"69",x"96",x"16",x"41",
x"67",x"54",x"04",x"80",x"90",x"81",x"C0",x"07",x"38",x"96",x"88",x"85",x"86",x"3F",
x"88",x"60",x"66",x"66",x"66",x"16",x"BF",x"56",x"20",x"07",x"33",x"33",x"83",x"3D",
x"31",x"82",x"32",x"08",x"84",x"19",x"BC",x"78",x"06",x"71",x"39",x"52",x"27",x"3A",
x"60",x"40",x"46",x"83",x"86",x"23",x"B8",x"00",x"00",x"00",x"07",x"36",x"22",x"3F",
x"00",x"00",x"00",x"27",x"44",x"89",x"3F",x"17",x"60",x"76",x"27",x"62",x"31",x"3F",
x"31",x"51",x"79",x"57",x"29",x"57",x"41",x"59",x"53",x"26",x"59",x"41",x"31",x"40",
x"79",x"26",x"63",x"79",x"70",x"15",x"40",x"20",x"51",x"75",x"19",x"47",x"10",x"40",
x"98",x"55",x"77",x"98",x"35",x"52",x"3F",x"00",x"00",x"00",x"80",x"76",x"32",x"44",
x"00",x"99",x"99",x"99",x"99",x"99",x"7E",x"F3",x"ED",x"56",x"3E",x"40",x"D3",x"02",
x"C3",x"33",x"02",x"3E",x"C0",x"D3",x"02",x"C3",x"3D",x"F1",x"3E",x"40",x"D3",x"02",
x"C3",x"41",x"C2",x"3E",x"50",x"D3",x"02",x"AF",x"01",x"60",x"04",x"ED",x"79",x"0C",
x"10",x"FB",x"21",x"45",x"C5",x"06",x"10",x"78",x"3D",x"D3",x"70",x"7E",x"D3",x"71",
x"23",x"10",x"F6",x"3E",x"80",x"D3",x"06",x"3A",x"22",x"0B",x"3C",x"20",x"04",x"32",
x"21",x"0B",x"3E",x"08",x"3C",x"28",x"4C",x"31",x"FF",x"BF",x"21",x"00",x"00",x"CD",
x"3E",x"C3",x"28",x"05",x"3D",x"D3",x"00",x"18",x"FB",x"31",x"AC",x"16",x"21",x"00",
x"80",x"CD",x"3E",x"C3",x"28",x"04",x"3E",x"88",x"ED",x"79",x"3E",x"70",x"D3",x"02",
x"21",x"00",x"40",x"CD",x"3E",x"C3",x"CC",x"3E",x"C3",x"2B",x"22",x"19",x"0B",x"3E",
x"40",x"D3",x"02",x"31",x"FF",x"BF",x"C3",x"A9",x"02",x"3E",x"80",x"D3",x"02",x"21",
x"00",x"C0",x"CD",x"38",x"03",x"3E",x"00",x"28",x"01",x"3D",x"08",x"18",x"07",x"67",
x"6F",x"2B",x"7C",x"B5",x"20",x"FB",x"3E",x"40",x"D3",x"02",x"C3",x"C9",x"02",x"3E",
x"C0",x"D3",x"02",x"31",x"AC",x"16",x"C3",x"00",x"F0",x"AF",x"32",x"11",x"0B",x"D3",
x"03",x"D3",x"07",x"D3",x"58",x"D3",x"59",x"D3",x"5A",x"D3",x"5B",x"D3",x"00",x"32",
x"4F",x"0B",x"3E",x"80",x"D3",x"06",x"32",x"13",x"0B",x"21",x"55",x"C5",x"01",x"70",
x"04",x"C5",x"5E",x"23",x"56",x"23",x"E5",x"EB",x"CD",x"21",x"C3",x"E1",x"C1",x"79",
x"D3",x"02",x"10",x"EF",x"3E",x"60",x"D3",x"02",x"C3",x"0D",x"03",x"3E",x"20",x"D3",
x"02",x"21",x"00",x"C0",x"11",x"34",x"03",x"06",x"04",x"1A",x"BE",x"20",x"05",x"13",
x"23",x"10",x"F8",x"E9",x"3E",x"60",x"D3",x"02",x"C3",x"29",x"C3",x"3E",x"70",x"D3",
x"02",x"32",x"03",x"00",x"FB",x"C3",x"EF",x"D9",x"4D",x"4F",x"50",x"53",x"E5",x"CD",
x"48",x"03",x"18",x"04",x"E5",x"CD",x"48",x"C3",x"D1",x"C0",x"EB",x"3E",x"AA",x"01",
x"3E",x"55",x"E5",x"5D",x"54",x"13",x"77",x"01",x"FF",x"3F",x"ED",x"B0",x"E1",x"06",
x"40",x"3D",x"35",x"ED",x"A1",x"2B",x"36",x"00",x"C0",x"23",x"E0",x"18",x"F5",x"E5",
x"DD",x"E5",x"FD",x"E5",x"D9",x"C5",x"D5",x"E5",x"D9",x"08",x"CD",x"7E",x"C3",x"D9",
x"E1",x"D1",x"C1",x"D9",x"FD",x"E1",x"DD",x"E1",x"E1",x"C3",x"37",x"0B",x"F5",x"C5",
x"D5",x"4F",x"B7",x"08",x"21",x"01",x"0B",x"7E",x"FE",x"02",x"20",x"01",x"35",x"11",
x"00",x"0B",x"79",x"07",x"38",x"03",x"11",x"08",x"0B",x"E6",x"E0",x"07",x"07",x"07",
x"47",x"79",x"E6",x"0F",x"4F",x"78",x"FE",x"07",x"28",x"32",x"68",x"AF",x"67",x"19",
x"3D",x"BE",x"20",x"05",x"79",x"FE",x"03",x"30",x"1D",x"7E",x"CB",x"BF",x"FE",x"07",
x"38",x"06",x"3E",x"FE",x"D1",x"C1",x"18",x"3C",x"CB",x"7E",x"28",x"06",x"21",x"66",
x"F1",x"C3",x"F0",x"FF",x"79",x"FE",x"03",x"30",x"01",x"46",x"78",x"FE",x"06",x"21",
x"6C",x"F1",x"28",x"EF",x"11",x"5D",x"C5",x"68",x"26",x"00",x"29",x"19",x"5E",x"23",
x"56",x"EB",x"7E",x"3D",x"B9",x"3E",x"FF",x"38",x"D1",x"23",x"EB",x"69",x"26",x"00",
x"29",x"19",x"5E",x"23",x"56",x"EB",x"08",x"D1",x"C1",x"CD",x"21",x"C3",x"B7",x"E1",
x"C8",x"F5",x"3A",x"20",x"0B",x"3C",x"28",x"0A",x"C5",x"D5",x"7C",x"21",x"E6",x"F1",
x"18",x"B9",x"D1",x"C1",x"F1",x"C9",x"3A",x"03",x"00",x"F5",x"E5",x"D5",x"C5",x"DD",
x"E5",x"FD",x"E5",x"08",x"F5",x"D9",x"E5",x"D5",x"C5",x"CD",x"37",x"C4",x"C1",x"D1",
x"E1",x"D9",x"F1",x"08",x"FD",x"E1",x"DD",x"E1",x"C1",x"D1",x"E1",x"F1",x"C3",x"41",
x"0B",x"3E",x"FF",x"32",x"20",x"0B",x"2A",x"1D",x"0B",x"23",x"22",x"1D",x"0B",x"3A",
x"4F",x"0B",x"D3",x"00",x"DB",x"59",x"4F",x"CB",x"67",x"CB",x"E1",x"D3",x"07",x"CC",
x"7D",x"C4",x"79",x"F6",x"F0",x"3C",x"28",x"1E",x"3A",x"1F",x"0B",x"0F",x"0F",x"61",
x"69",x"01",x"58",x"04",x"57",x"AF",x"CB",x"0A",x"1F",x"CB",x"0C",x"38",x"02",x"ED",
x"79",x"0C",x"10",x"F3",x"4D",x"21",x"78",x"C4",x"18",x"2B",x"AF",x"32",x"20",x"0B",
x"C9",x"C5",x"3A",x"10",x"0B",x"4F",x"06",x"04",x"CB",x"19",x"C5",x"38",x"10",x"3E",
x"04",x"90",x"47",x"0E",x"00",x"21",x"99",x"C4",x"E5",x"E5",x"E5",x"E5",x"C3",x"D8",
x"C3",x"3E",x"70",x"D3",x"02",x"C1",x"10",x"E4",x"21",x"AA",x"C4",x"E5",x"21",x"27",
x"F2",x"C3",x"F0",x"FF",x"C1",x"C9",x"05",x"09",x"C5",x"B7",x"C4",x"D0",x"C4",x"E2",
x"C4",x"0E",x"C5",x"2A",x"19",x"0B",x"3E",x"FB",x"B7",x"ED",x"52",x"D8",x"E5",x"11",
x"AC",x"1E",x"ED",x"52",x"E1",x"D8",x"54",x"5D",x"13",x"22",x"19",x"0B",x"AF",x"C9",
x"21",x"07",x"0B",x"04",x"28",x"03",x"21",x"0F",x"0B",x"E5",x"CD",x"0E",x"C5",x"E1",
x"B7",x"C0",x"71",x"C9",x"21",x"00",x"0B",x"14",x"28",x"03",x"21",x"08",x"0B",x"E5",
x"3E",x"06",x"B8",x"38",x"19",x"58",x"16",x"00",x"19",x"5E",x"1C",x"28",x"11",x"D1",
x"E5",x"EB",x"B9",x"38",x"0B",x"59",x"AF",x"57",x"19",x"5E",x"1C",x"28",x"03",x"E1",
x"71",x"C9",x"E1",x"3E",x"FE",x"C9",x"D5",x"DD",x"21",x"40",x"00",x"06",x"04",x"DD",
x"E5",x"E1",x"C5",x"1A",x"3C",x"47",x"1A",x"BE",x"20",x"17",x"23",x"13",x"10",x"F8",
x"C1",x"DD",x"E5",x"E1",x"11",x"07",x"00",x"19",x"7E",x"B9",x"20",x"08",x"3E",x"04",
x"90",x"4F",x"AF",x"D1",x"C9",x"C1",x"11",x"30",x"00",x"DD",x"19",x"D1",x"D5",x"10",
x"D4",x"3E",x"FD",x"18",x"F0",x"FF",x"0E",x"00",x"00",x"03",x"03",x"03",x"00",x"42",
x"3C",x"02",x"4D",x"32",x"4B",x"40",x"63",x"F2",x"C9",x"EC",x"D5",x"60",x"D9",x"E2",
x"D9",x"74",x"C9",x"E3",x"D5",x"98",x"CF",x"2A",x"D9",x"FF",x"D8",x"BB",x"D9",x"00",
x"00",x"AC",x"C4",x"EB",x"E5",x"D5",x"C5",x"E5",x"D5",x"EB",x"2A",x"19",x"0B",x"B7",
x"ED",x"52",x"3E",x"FA",x"D1",x"E1",x"D8",x"4E",x"EB",x"CD",x"8E",x"C5",x"C1",x"D1",
x"E1",x"B7",x"C0",x"ED",x"A1",x"E0",x"18",x"E0",x"E9",x"E5",x"D5",x"C5",x"E5",x"D5",
x"2A",x"19",x"0B",x"B7",x"ED",x"52",x"3E",x"FA",x"D1",x"E1",x"D8",x"CD",x"8E",x"C5",
x"08",x"79",x"C1",x"D1",x"E1",x"08",x"B7",x"C0",x"08",x"12",x"AF",x"EB",x"ED",x"A1",
x"EB",x"E0",x"18",x"DB",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"18",x"18",x"18",x"18",x"18",x"00",x"18",x"00",x"00",x"00",x"36",x"36",x"36",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"36",x"7F",x"36",x"7F",x"36",x"36",
x"00",x"00",x"00",x"18",x"3E",x"58",x"3C",x"1A",x"7C",x"18",x"00",x"00",x"00",x"60",
x"66",x"0C",x"18",x"30",x"66",x"06",x"00",x"00",x"00",x"10",x"28",x"28",x"30",x"54",
x"48",x"34",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"0C",x"18",x"30",x"30",x"30",x"18",x"0C",x"00",x"00",x"00",x"30",x"18",x"0C",
x"0C",x"0C",x"18",x"30",x"00",x"00",x"00",x"00",x"10",x"54",x"38",x"38",x"54",x"10",
x"00",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"18",x"18",x"30",x"00",x"00",x"00",x"00",x"00",x"7C",x"7C",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",
x"00",x"00",x"06",x"0C",x"18",x"30",x"60",x"00",x"00",x"00",x"00",x"3C",x"66",x"6E",
x"7E",x"76",x"66",x"3C",x"00",x"00",x"00",x"18",x"38",x"18",x"18",x"18",x"18",x"18",
x"00",x"00",x"00",x"3C",x"66",x"06",x"1C",x"30",x"60",x"7E",x"00",x"00",x"00",x"7E",
x"06",x"0C",x"1C",x"06",x"46",x"3C",x"00",x"00",x"00",x"0C",x"1C",x"2C",x"4C",x"7E",
x"0C",x"0C",x"00",x"00",x"00",x"7E",x"60",x"7C",x"06",x"06",x"46",x"3C",x"00",x"00",
x"00",x"3C",x"60",x"60",x"7C",x"66",x"66",x"3C",x"00",x"00",x"00",x"7E",x"06",x"0C",
x"18",x"30",x"60",x"60",x"00",x"00",x"00",x"3C",x"66",x"66",x"3C",x"66",x"66",x"3C",
x"00",x"00",x"00",x"3C",x"66",x"66",x"3E",x"06",x"0C",x"38",x"00",x"00",x"00",x"00",
x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",
x"18",x"18",x"30",x"00",x"00",x"06",x"0C",x"18",x"30",x"18",x"0C",x"06",x"00",x"00",
x"00",x"00",x"00",x"7C",x"00",x"7C",x"00",x"00",x"00",x"00",x"00",x"30",x"18",x"0C",
x"06",x"0C",x"18",x"30",x"00",x"00",x"00",x"3C",x"66",x"06",x"0C",x"18",x"00",x"18",
x"00",x"00",x"00",x"3E",x"63",x"67",x"6B",x"6F",x"60",x"3C",x"00",x"00",x"00",x"1C",
x"3E",x"63",x"63",x"7F",x"63",x"63",x"00",x"00",x"00",x"7E",x"63",x"63",x"7E",x"63",
x"63",x"7E",x"00",x"00",x"00",x"3E",x"63",x"60",x"60",x"60",x"63",x"3E",x"00",x"00",
x"00",x"7E",x"33",x"33",x"33",x"33",x"33",x"7E",x"00",x"00",x"00",x"7E",x"60",x"60",
x"7C",x"60",x"60",x"7E",x"00",x"00",x"00",x"7E",x"60",x"60",x"7C",x"60",x"60",x"60",
x"00",x"00",x"00",x"3E",x"63",x"60",x"60",x"67",x"63",x"3E",x"00",x"00",x"00",x"63",
x"63",x"63",x"7F",x"63",x"63",x"63",x"00",x"00",x"00",x"3C",x"18",x"18",x"18",x"18",
x"18",x"3C",x"00",x"00",x"00",x"06",x"06",x"06",x"06",x"66",x"66",x"3C",x"00",x"00",
x"00",x"63",x"66",x"6C",x"78",x"6C",x"66",x"63",x"00",x"00",x"00",x"60",x"60",x"60",
x"60",x"60",x"60",x"7E",x"00",x"00",x"00",x"63",x"77",x"6B",x"63",x"63",x"63",x"63",
x"00",x"00",x"00",x"66",x"66",x"76",x"6E",x"66",x"66",x"66",x"00",x"00",x"00",x"3E",
x"63",x"63",x"63",x"63",x"63",x"3E",x"00",x"00",x"00",x"7E",x"63",x"63",x"7E",x"60",
x"60",x"60",x"00",x"00",x"00",x"3E",x"63",x"63",x"63",x"6B",x"67",x"3E",x"01",x"00",
x"00",x"7E",x"63",x"63",x"7E",x"6C",x"66",x"63",x"00",x"00",x"00",x"3E",x"63",x"60",
x"3E",x"03",x"63",x"3E",x"00",x"00",x"00",x"7E",x"5A",x"18",x"18",x"18",x"18",x"18",
x"00",x"00",x"00",x"63",x"63",x"63",x"63",x"63",x"63",x"3E",x"00",x"00",x"00",x"63",
x"63",x"63",x"63",x"36",x"1C",x"08",x"00",x"00",x"00",x"63",x"63",x"63",x"6B",x"6B",
x"3E",x"14",x"00",x"00",x"00",x"66",x"66",x"3C",x"18",x"3C",x"66",x"66",x"00",x"00",
x"00",x"66",x"66",x"3C",x"18",x"18",x"18",x"18",x"00",x"00",x"00",x"7E",x"06",x"0C",
x"18",x"30",x"60",x"7E",x"00",x"00",x"00",x"3C",x"30",x"30",x"30",x"30",x"30",x"3C",
x"00",x"00",x"00",x"00",x"60",x"30",x"18",x"0C",x"06",x"00",x"00",x"00",x"00",x"3C",
x"0C",x"0C",x"0C",x"0C",x"0C",x"3C",x"00",x"00",x"00",x"18",x"3C",x"66",x"42",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"00",x"00",
x"00",x"30",x"30",x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",
x"06",x"3E",x"66",x"3E",x"00",x"00",x"00",x"60",x"60",x"7C",x"66",x"66",x"66",x"7C",
x"00",x"00",x"00",x"00",x"00",x"1E",x"30",x"30",x"30",x"1E",x"00",x"00",x"00",x"06",
x"06",x"3E",x"66",x"66",x"66",x"3E",x"00",x"00",x"00",x"00",x"00",x"3C",x"66",x"7E",
x"60",x"3C",x"00",x"00",x"00",x"0C",x"18",x"18",x"3C",x"18",x"18",x"18",x"00",x"00",
x"00",x"00",x"00",x"3E",x"66",x"66",x"66",x"3E",x"06",x"3C",x"00",x"60",x"60",x"7C",
x"66",x"66",x"66",x"66",x"00",x"00",x"00",x"18",x"00",x"38",x"18",x"18",x"18",x"3C",
x"00",x"00",x"00",x"18",x"00",x"38",x"18",x"18",x"18",x"18",x"18",x"70",x"00",x"60",
x"60",x"66",x"6C",x"78",x"6C",x"66",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",
x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"76",x"6B",x"6B",x"6B",x"6B",x"00",x"00",
x"00",x"00",x"00",x"7C",x"66",x"66",x"66",x"66",x"00",x"00",x"00",x"00",x"00",x"3C",
x"66",x"66",x"66",x"3C",x"00",x"00",x"00",x"00",x"00",x"7C",x"66",x"66",x"66",x"7C",
x"60",x"60",x"00",x"00",x"00",x"3E",x"66",x"66",x"66",x"3E",x"06",x"06",x"00",x"00",
x"00",x"36",x"38",x"30",x"30",x"30",x"00",x"00",x"00",x"00",x"00",x"1E",x"30",x"1C",
x"06",x"3C",x"00",x"00",x"00",x"18",x"18",x"3C",x"18",x"18",x"18",x"0C",x"00",x"00",
x"00",x"00",x"00",x"66",x"66",x"66",x"66",x"3E",x"00",x"00",x"00",x"00",x"00",x"66",
x"66",x"66",x"3C",x"18",x"00",x"00",x"00",x"00",x"00",x"63",x"63",x"6B",x"3E",x"14",
x"00",x"00",x"00",x"00",x"00",x"66",x"3C",x"18",x"3C",x"66",x"00",x"00",x"00",x"00",
x"00",x"66",x"66",x"66",x"66",x"3E",x"06",x"3C",x"00",x"00",x"00",x"7E",x"0C",x"18",
x"30",x"7E",x"00",x"00",x"00",x"0E",x"18",x"18",x"70",x"18",x"18",x"0E",x"00",x"00",
x"00",x"18",x"18",x"18",x"00",x"18",x"18",x"18",x"00",x"00",x"00",x"70",x"18",x"18",
x"0E",x"18",x"18",x"70",x"00",x"00",x"00",x"00",x"00",x"33",x"6B",x"66",x"00",x"00",
x"00",x"00",x"00",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"0D",x"A9",
x"C9",x"94",x"CC",x"86",x"CC",x"4B",x"CF",x"F4",x"C9",x"49",x"CA",x"DA",x"CA",x"D7",
x"CA",x"F3",x"CB",x"FF",x"CB",x"48",x"CD",x"2C",x"CF",x"38",x"CA",x"E1",x"3A",x"03",
x"00",x"F5",x"3E",x"50",x"32",x"03",x"00",x"D3",x"02",x"E5",x"21",x"A1",x"C9",x"E3",
x"E9",x"08",x"F1",x"32",x"03",x"00",x"D3",x"02",x"08",x"C9",x"87",x"5F",x"16",x"00",
x"19",x"5E",x"23",x"56",x"C9",x"21",x"FF",x"03",x"B7",x"ED",x"42",x"C9",x"21",x"BF",
x"03",x"B7",x"ED",x"52",x"C9",x"3A",x"73",x"0B",x"47",x"04",x"CB",x"3C",x"CB",x"1D",
x"10",x"FA",x"C9",x"CD",x"6D",x"CB",x"CD",x"05",x"CC",x"32",x"93",x"0B",x"11",x"40",
x"00",x"CD",x"8F",x"CB",x"CD",x"0D",x"CC",x"32",x"94",x"0B",x"3A",x"75",x"0B",x"4F",
x"2A",x"76",x"0B",x"C9",x"00",x"50",x"44",x"41",x"00",x"55",x"50",x"44",x"0E",x"01",
x"79",x"FE",x"03",x"3E",x"F7",x"D0",x"AF",x"32",x"4B",x"0B",x"32",x"4E",x"0B",x"32",
x"50",x"0B",x"3C",x"32",x"4C",x"0B",x"B9",x"30",x"0A",x"DB",x"59",x"07",x"07",x"3E",
x"0F",x"30",x"02",x"3E",x"0C",x"32",x"4D",x"0B",x"79",x"32",x"73",x"0B",x"C5",x"CD",
x"49",x"CA",x"C1",x"79",x"21",x"13",x"0B",x"AE",x"E6",x"FC",x"A9",x"77",x"D3",x"06",
x"DB",x"59",x"07",x"07",x"11",x"EE",x"C9",x"30",x"03",x"11",x"EA",x"C9",x"1A",x"D3",
x"60",x"13",x"1A",x"D3",x"61",x"13",x"1A",x"D3",x"62",x"13",x"1A",x"D3",x"63",x"AF",
x"C9",x"CD",x"8F",x"C9",x"CD",x"D4",x"CF",x"CD",x"05",x"CC",x"21",x"00",x"80",x"11",
x"01",x"80",x"77",x"01",x"FF",x"3B",x"ED",x"B0",x"CD",x"FF",x"CB",x"47",x"4F",x"57",
x"5F",x"ED",x"53",x"7E",x"0B",x"ED",x"43",x"7C",x"0B",x"2A",x"7C",x"0B",x"E5",x"06",
x"04",x"CD",x"C6",x"C9",x"E3",x"CD",x"C1",x"C9",x"22",x"78",x"0B",x"4F",x"7D",x"21",
x"B4",x"CA",x"09",x"E6",x"07",x"3C",x"47",x"7E",x"1E",x"0F",x"10",x"FD",x"32",x"75",
x"0B",x"ED",x"5B",x"7E",x"0B",x"21",x"BF",x"03",x"AF",x"ED",x"52",x"06",x"02",x"CD",
x"C6",x"C9",x"22",x"7A",x"0B",x"65",x"CB",x"3C",x"1F",x"CB",x"3C",x"1F",x"6F",x"C1",
x"09",x"11",x"00",x"80",x"19",x"22",x"76",x"0B",x"AF",x"C9",x"80",x"88",x"AA",x"30",
x"0C",x"E6",x"01",x"28",x"03",x"C9",x"30",x"08",x"3A",x"94",x"0B",x"FD",x"E9",x"E6",
x"02",x"C0",x"3A",x"93",x"0B",x"FD",x"E9",x"A6",x"AE",x"A1",x"AE",x"77",x"C9",x"A1",
x"B6",x"77",x"C9",x"CD",x"7A",x"CC",x"CD",x"8F",x"C9",x"3E",x"F9",x"CD",x"B3",x"C9",
x"D4",x"BA",x"C9",x"D8",x"3A",x"74",x"0B",x"B7",x"CA",x"65",x"CA",x"D9",x"ED",x"4B",
x"78",x"0B",x"ED",x"5B",x"7A",x"0B",x"C5",x"D5",x"CD",x"CD",x"C9",x"D9",x"CD",x"65",
x"CA",x"ED",x"4B",x"78",x"0B",x"ED",x"5B",x"7A",x"0B",x"AF",x"EB",x"D1",x"CD",x"61",
x"CB",x"D1",x"E5",x"60",x"69",x"CD",x"61",x"CB",x"E5",x"21",x"DB",x"CB",x"CD",x"AA",
x"C9",x"ED",x"53",x"86",x"0B",x"E1",x"D1",x"E5",x"ED",x"52",x"E1",x"38",x"01",x"EB",
x"44",x"4D",x"D5",x"CE",x"00",x"ED",x"52",x"E5",x"CB",x"3A",x"CB",x"1B",x"19",x"E5",
x"21",x"E3",x"CB",x"CD",x"AA",x"C9",x"ED",x"53",x"84",x"0B",x"E1",x"D1",x"D9",x"E3",
x"7C",x"45",x"04",x"3C",x"08",x"E1",x"18",x"04",x"08",x"CD",x"A8",x"CB",x"3A",x"83",
x"0B",x"07",x"32",x"83",x"0B",x"CD",x"BE",x"CA",x"10",x"F1",x"08",x"3D",x"20",x"EC",
x"C9",x"ED",x"52",x"30",x"06",x"EB",x"21",x"01",x"00",x"ED",x"52",x"17",x"C9",x"3A",
x"4C",x"0B",x"3D",x"E6",x"0F",x"4F",x"21",x"7F",x"CB",x"06",x"00",x"09",x"7E",x"32",
x"83",x"0B",x"C9",x"FF",x"AA",x"CC",x"EE",x"88",x"DA",x"E4",x"F6",x"FA",x"FE",x"FC",
x"F8",x"F0",x"EA",x"FF",x"FF",x"D5",x"3A",x"4B",x"0B",x"E6",x"03",x"21",x"A0",x"CB",
x"CD",x"AA",x"C9",x"D5",x"FD",x"E1",x"D1",x"C9",x"CE",x"CA",x"D3",x"CA",x"CD",x"CA",
x"CF",x"CA",x"D9",x"CB",x"7C",x"28",x"08",x"09",x"D9",x"DD",x"2A",x"84",x"0B",x"DD",
x"E9",x"19",x"D9",x"DD",x"2A",x"86",x"0B",x"DD",x"E9",x"B7",x"ED",x"52",x"CB",x"01",
x"D0",x"2D",x"C9",x"CB",x"09",x"30",x"01",x"2C",x"B7",x"ED",x"52",x"C9",x"CB",x"01",
x"30",x"01",x"2D",x"19",x"C9",x"19",x"CB",x"09",x"D0",x"2C",x"C9",x"D5",x"CB",x"CE",
x"CB",x"C5",x"CB",x"BD",x"CB",x"D6",x"CB",x"D3",x"CB",x"C0",x"CB",x"D3",x"CB",x"D6",
x"CB",x"CA",x"CB",x"C0",x"CB",x"CA",x"CB",x"CD",x"8F",x"C9",x"CD",x"D9",x"C9",x"CD",
x"C0",x"CA",x"3E",x"FF",x"26",x"AF",x"32",x"74",x"0B",x"AF",x"C9",x"3A",x"4E",x"0B",
x"CD",x"10",x"CC",x"47",x"C9",x"3A",x"4D",x"0B",x"2A",x"73",x"0B",x"CB",x"3D",x"38",
x"09",x"CB",x"3D",x"38",x"16",x"E6",x"01",x"1F",x"9F",x"C9",x"E6",x"03",x"1F",x"CB",
x"15",x"1F",x"9F",x"CB",x"1D",x"1F",x"CB",x"2F",x"CB",x"2F",x"CB",x"2F",x"C9",x"E6",
x"0F",x"26",x"04",x"1F",x"CB",x"1D",x"CB",x"2D",x"25",x"20",x"F8",x"7D",x"C9",x"CD",
x"E2",x"C9",x"3A",x"73",x"0B",x"47",x"79",x"A6",x"CB",x"38",x"38",x"0A",x"CB",x"38",
x"38",x"15",x"C6",x"FF",x"17",x"E6",x"01",x"C9",x"C6",x"F0",x"CB",x"11",x"E6",x"0F",
x"C6",x"FF",x"17",x"CB",x"19",x"17",x"E6",x"03",x"C9",x"C6",x"C0",x"17",x"E6",x"7F",
x"C6",x"E0",x"17",x"E6",x"3F",x"C6",x"F0",x"17",x"E6",x"1F",x"C6",x"F8",x"17",x"E6",
x"0F",x"C9",x"2A",x"7C",x"0B",x"09",x"44",x"4D",x"2A",x"7E",x"0B",x"19",x"EB",x"C9",
x"EB",x"E5",x"C5",x"4E",x"CD",x"94",x"CC",x"C1",x"E1",x"ED",x"A1",x"E0",x"18",x"F3",
x"CD",x"8F",x"C9",x"79",x"FE",x"20",x"30",x"0C",x"FE",x"0A",x"CA",x"31",x"CD",x"FE",
x"0D",x"CA",x"2B",x"CD",x"AF",x"C9",x"FE",x"E0",x"3E",x"00",x"D0",x"D9",x"11",x"DC",
x"FF",x"3A",x"73",x"0B",x"47",x"3E",x"01",x"04",x"87",x"10",x"FD",x"32",x"82",x"0B",
x"6F",x"87",x"85",x"87",x"85",x"4F",x"AF",x"CD",x"7A",x"CC",x"CD",x"BA",x"C9",x"D8",
x"CD",x"B3",x"C9",x"30",x"06",x"CD",x"2B",x"CD",x"CD",x"31",x"CD",x"CD",x"D0",x"C9",
x"D9",x"11",x"74",x"C4",x"CB",x"79",x"28",x"03",x"11",x"40",x"07",x"CB",x"B9",x"06",
x"00",x"60",x"69",x"29",x"29",x"09",x"29",x"19",x"06",x"0A",x"3A",x"50",x"0B",x"5F",
x"2B",x"23",x"4E",x"D9",x"06",x"08",x"18",x"03",x"CD",x"D6",x"CB",x"D9",x"CB",x"11",
x"7B",x"D9",x"CD",x"B7",x"CA",x"10",x"F3",x"CD",x"D3",x"CB",x"06",x"07",x"CD",x"C0",
x"CB",x"10",x"FB",x"D9",x"10",x"DF",x"3A",x"82",x"0B",x"87",x"87",x"87",x"4F",x"CD",
x"7A",x"CC",x"CD",x"B3",x"C9",x"30",x"07",x"01",x"31",x"CD",x"C5",x"01",x"00",x"00",
x"C3",x"69",x"CA",x"11",x"B4",x"FF",x"CD",x"7A",x"CC",x"AF",x"CD",x"BA",x"C9",x"D8",
x"11",x"D8",x"FF",x"01",x"00",x"00",x"CD",x"7A",x"CC",x"C3",x"65",x"CA",x"CD",x"8F",
x"C9",x"ED",x"73",x"88",x"0B",x"FD",x"21",x"CF",x"CA",x"CD",x"3F",x"CC",x"CD",x"10",
x"CC",x"32",x"8A",x"0B",x"5F",x"CD",x"0D",x"CC",x"AB",x"21",x"00",x"00",x"C8",x"22",
x"91",x"0B",x"E5",x"2A",x"7C",x"0B",x"06",x"04",x"CD",x"C6",x"C9",x"E5",x"CD",x"DF",
x"C9",x"3E",x"40",x"D1",x"93",x"47",x"22",x"8D",x"0B",x"ED",x"43",x"8B",x"0B",x"06",
x"01",x"18",x"1E",x"E1",x"7C",x"B5",x"C8",x"C1",x"22",x"91",x"0B",x"ED",x"43",x"8B",
x"0B",x"E1",x"11",x"40",x"00",x"19",x"22",x"8D",x"0B",x"06",x"02",x"11",x"00",x"BC",
x"ED",x"52",x"D2",x"63",x"CE",x"D9",x"CD",x"92",x"CE",x"38",x"DC",x"2A",x"91",x"0B",
x"7C",x"CB",x"BC",x"CB",x"B4",x"22",x"8F",x"0B",x"EB",x"CB",x"77",x"28",x"09",x"07",
x"D9",x"A8",x"D9",x"E6",x"01",x"C2",x"62",x"CE",x"2A",x"8D",x"0B",x"ED",x"4B",x"8B",
x"0B",x"3A",x"8A",x"0B",x"AE",x"A1",x"20",x"5F",x"3E",x"40",x"90",x"3C",x"47",x"11",
x"00",x"00",x"18",x"0B",x"3A",x"8A",x"0B",x"AE",x"A1",x"20",x"0B",x"CD",x"C0",x"CA",
x"13",x"CB",x"01",x"30",x"F1",x"2D",x"10",x"EE",x"3E",x"40",x"90",x"3C",x"47",x"CB",
x"09",x"30",x"02",x"2C",x"05",x"E5",x"C5",x"D5",x"2A",x"8D",x"0B",x"ED",x"4B",x"8B",
x"0B",x"CD",x"7A",x"CE",x"E3",x"7C",x"B5",x"28",x"02",x"CB",x"FC",x"19",x"E3",x"E5",
x"2A",x"8F",x"0B",x"B7",x"ED",x"52",x"D1",x"E3",x"F5",x"3E",x"80",x"CB",x"7C",x"20",
x"09",x"38",x"09",x"D9",x"CB",x"08",x"CB",x"00",x"D9",x"1F",x"AC",x"67",x"F1",x"E3",
x"38",x"36",x"28",x"34",x"EB",x"CD",x"92",x"CE",x"DA",x"85",x"CD",x"7B",x"B7",x"20",
x"01",x"15",x"3A",x"8A",x"0B",x"AE",x"A1",x"28",x"0B",x"1D",x"28",x"1A",x"CB",x"09",
x"30",x"F2",x"2C",x"05",x"18",x"EE",x"7B",x"B7",x"20",x"01",x"14",x"ED",x"53",x"8F",
x"0B",x"E5",x"E3",x"C5",x"CD",x"7A",x"CE",x"D5",x"18",x"AF",x"15",x"F2",x"44",x"CE",
x"D9",x"05",x"CA",x"85",x"CD",x"D9",x"2A",x"8D",x"0B",x"11",x"80",x"FF",x"19",x"22",
x"8D",x"0B",x"CB",x"7C",x"CA",x"85",x"CD",x"C3",x"A4",x"CD",x"11",x"00",x"00",x"3A",
x"8A",x"0B",x"AE",x"A1",x"C0",x"13",x"3A",x"94",x"0B",x"A1",x"AE",x"77",x"CB",x"09",
x"30",x"EF",x"2C",x"10",x"EC",x"C9",x"E5",x"D5",x"21",x"EA",x"FF",x"39",x"ED",x"5B",
x"17",x"0B",x"ED",x"52",x"D2",x"C9",x"CE",x"C5",x"D9",x"C5",x"2A",x"88",x"0B",x"2B",
x"2B",x"2B",x"54",x"5D",x"4D",x"44",x"21",x"09",x"00",x"39",x"B7",x"ED",x"42",x"60",
x"69",x"20",x"13",x"01",x"0A",x"00",x"ED",x"B8",x"EB",x"F9",x"33",x"B7",x"EB",x"ED",
x"52",x"3F",x"C1",x"D9",x"C1",x"D1",x"E1",x"C9",x"CD",x"FE",x"CE",x"09",x"01",x"00",
x"BC",x"ED",x"42",x"30",x"06",x"09",x"CD",x"14",x"CF",x"28",x"0F",x"CD",x"FD",x"CE",
x"B7",x"ED",x"42",x"01",x"00",x"80",x"ED",x"42",x"09",x"D4",x"14",x"CF",x"D9",x"01",
x"06",x"00",x"20",x"05",x"ED",x"B8",x"C3",x"AC",x"CE",x"B7",x"ED",x"42",x"C3",x"AC",
x"CE",x"D9",x"E5",x"D9",x"E1",x"56",x"2B",x"5E",x"2B",x"2B",x"46",x"2B",x"7E",x"E6",
x"3F",x"2B",x"6E",x"67",x"78",x"01",x"40",x"00",x"EB",x"C9",x"4F",x"3A",x"8A",x"0B",
x"47",x"78",x"AE",x"A1",x"C8",x"1D",x"28",x"07",x"CB",x"09",x"30",x"F5",x"23",x"18",
x"F2",x"15",x"F2",x"20",x"CF",x"C9",x"79",x"FE",x"E0",x"30",x"01",x"B7",x"3E",x"F8",
x"F0",x"CB",x"B9",x"06",x"00",x"69",x"60",x"29",x"29",x"09",x"29",x"01",x"40",x"07",
x"09",x"EB",x"01",x"0A",x"00",x"ED",x"B0",x"AF",x"C9",x"C5",x"21",x"00",x"00",x"05",
x"FA",x"54",x"CF",x"68",x"3A",x"73",x"0B",x"C6",x"04",x"47",x"29",x"10",x"FD",x"E5",
x"11",x"D8",x"FF",x"21",x"BF",x"03",x"41",x"05",x"FA",x"6E",x"CF",x"28",x"03",x"19",
x"10",x"FD",x"EB",x"C1",x"D9",x"ED",x"4B",x"7C",x"0B",x"ED",x"5B",x"7E",x"0B",x"D9",
x"E1",x"7D",x"B7",x"20",x"04",x"D9",x"D5",x"D9",x"D1",x"7C",x"B7",x"20",x"04",x"D9",
x"C5",x"D9",x"C1",x"3E",x"F9",x"CD",x"B3",x"C9",x"D8",x"CD",x"BA",x"C9",x"D8",x"C3",
x"65",x"CA",x"05",x"A3",x"CF",x"52",x"D0",x"41",x"D0",x"1D",x"D0",x"13",x"D0",x"3E",
x"50",x"D3",x"02",x"21",x"48",x"0E",x"ED",x"4B",x"49",x"0E",x"34",x"3E",x"94",x"96",
x"28",x"1C",x"FE",x"80",x"C0",x"77",x"3A",x"66",x"0B",x"16",x"7F",x"B7",x"28",x"0C",
x"16",x"9E",x"0F",x"38",x"07",x"16",x"9F",x"0F",x"38",x"02",x"16",x"8F",x"7A",x"C3",
x"20",x"D4",x"77",x"C3",x"91",x"D4",x"21",x"48",x"0E",x"06",x"20",x"AF",x"77",x"23",
x"10",x"FC",x"21",x"01",x"01",x"22",x"49",x"0E",x"21",x"00",x"01",x"11",x"01",x"01",
x"01",x"FF",x"05",x"36",x"20",x"ED",x"B0",x"3A",x"73",x"0B",x"87",x"87",x"21",x"07",
x"D0",x"4F",x"09",x"11",x"68",x"0E",x"3E",x"C3",x"12",x"13",x"0E",x"04",x"ED",x"B0",
x"C9",x"AD",x"D3",x"40",x"01",x"BC",x"D3",x"20",x"02",x"D9",x"D3",x"10",x"04",x"2A",
x"49",x"0E",x"22",x"4E",x"0E",x"3E",x"80",x"18",x"1C",x"2A",x"49",x"0E",x"78",x"B7",
x"28",x"07",x"3A",x"6B",x"0E",x"B8",x"38",x"14",x"60",x"79",x"B7",x"28",x"06",x"3E",
x"18",x"B9",x"38",x"0A",x"69",x"22",x"49",x"0E",x"AF",x"32",x"4D",x"0E",x"AF",x"C9",
x"3E",x"F6",x"C9",x"D9",x"CD",x"49",x"D4",x"D9",x"21",x"B7",x"D0",x"F2",x"6D",x"C5",
x"21",x"58",x"D0",x"C3",x"8F",x"C5",x"CD",x"49",x"D4",x"F2",x"B7",x"D0",x"3E",x"50",
x"32",x"03",x"00",x"D3",x"02",x"3A",x"4D",x"0E",x"0F",x"DA",x"FA",x"D0",x"CD",x"9C",
x"D3",x"ED",x"4B",x"49",x"0E",x"C5",x"ED",x"5B",x"4E",x"0E",x"79",x"BB",x"38",x"06",
x"20",x"09",x"78",x"BA",x"30",x"0F",x"CD",x"38",x"D0",x"18",x"0A",x"0D",x"28",x"F8",
x"2B",x"CB",x"7E",x"16",x"01",x"20",x"E7",x"C1",x"CD",x"77",x"D4",x"3E",x"13",x"32",
x"48",x"0E",x"21",x"10",x"0B",x"CB",x"96",x"F7",x"91",x"CB",x"D6",x"F5",x"C5",x"ED",
x"4B",x"49",x"0E",x"CD",x"91",x"D4",x"C1",x"F1",x"C0",x"79",x"FE",x"1B",x"28",x"8A",
x"FE",x"0D",x"28",x"39",x"CD",x"24",x"D1",x"18",x"AF",x"3E",x"50",x"32",x"03",x"00",
x"D3",x"02",x"21",x"38",x"D0",x"E5",x"79",x"FE",x"0D",x"20",x"06",x"3E",x"01",x"32",
x"4A",x"0E",x"C9",x"FE",x"0A",x"20",x"15",x"ED",x"4B",x"49",x"0E",x"79",x"CD",x"9F",
x"D3",x"0C",x"38",x"F9",x"0D",x"C5",x"CD",x"63",x"D3",x"F1",x"32",x"4A",x"0E",x"C9",
x"CD",x"24",x"D1",x"AF",x"C9",x"3A",x"4D",x"0E",x"07",x"ED",x"4B",x"4E",x"0E",x"D4",
x"70",x"D3",x"ED",x"43",x"49",x"0E",x"ED",x"4B",x"49",x"0E",x"79",x"CD",x"9F",x"D3",
x"B8",x"38",x"17",x"CD",x"84",x"D3",x"04",x"3A",x"6B",x"0E",x"B8",x"30",x"03",x"06",
x"01",x"0C",x"ED",x"43",x"49",x"0E",x"4E",x"3E",x"01",x"C3",x"39",x"D0",x"CD",x"63",
x"D3",x"0E",x"0D",x"C3",x"38",x"D0",x"FE",x"20",x"38",x"2F",x"FE",x"E0",x"30",x"2B",
x"08",x"CD",x"84",x"D3",x"08",x"77",x"ED",x"4B",x"49",x"0E",x"C5",x"CD",x"20",x"D4",
x"C1",x"79",x"CD",x"9F",x"D3",x"B8",x"30",x"01",x"70",x"04",x"3A",x"6B",x"0E",x"B8",
x"30",x"08",x"06",x"01",x"0C",x"CB",x"7E",x"CC",x"CB",x"D2",x"ED",x"43",x"49",x"0E",
x"C9",x"21",x"70",x"D1",x"06",x"0B",x"BE",x"23",x"5E",x"23",x"56",x"23",x"28",x"03",
x"10",x"F6",x"C9",x"ED",x"4B",x"49",x"0E",x"3A",x"6B",x"0E",x"EB",x"E9",x"13",x"91",
x"D1",x"04",x"98",x"D1",x"05",x"95",x"D1",x"18",x"9E",x"D1",x"16",x"05",x"D2",x"07",
x"87",x"D2",x"08",x"78",x"D2",x"19",x"FD",x"D1",x"0E",x"F7",x"D1",x"0B",x"A8",x"D1",
x"09",x"CD",x"D1",x"05",x"20",x"0F",x"47",x"0D",x"18",x"0A",x"04",x"B8",x"30",x"07",
x"06",x"01",x"0C",x"79",x"FE",x"19",x"C8",x"ED",x"43",x"49",x"0E",x"C9",x"C5",x"CD",
x"AD",x"D4",x"C1",x"CD",x"84",x"D3",x"05",x"3A",x"6B",x"0E",x"90",x"36",x"20",x"23",
x"3D",x"20",x"FA",x"CD",x"9C",x"D3",x"70",x"0C",x"23",x"D0",x"46",x"79",x"D9",x"CD",
x"1E",x"D3",x"D9",x"CB",x"00",x"18",x"F4",x"CD",x"9C",x"D3",x"08",x"78",x"3D",x"E6",
x"F8",x"C6",x"09",x"47",x"3A",x"6B",x"0E",x"B8",x"30",x"0A",x"F6",x"80",x"77",x"06",
x"01",x"0C",x"08",x"D4",x"CB",x"D2",x"79",x"CD",x"9F",x"D3",x"05",x"B8",x"30",x"01",
x"70",x"04",x"ED",x"43",x"49",x"0E",x"C9",x"CD",x"70",x"D3",x"C3",x"D6",x"D2",x"CD",
x"70",x"D3",x"CD",x"9C",x"D3",x"18",x"BD",x"CD",x"9C",x"D3",x"B8",x"D8",x"1E",x"01",
x"18",x"02",x"23",x"1C",x"7E",x"07",x"0C",x"38",x"F9",x"34",x"3A",x"6B",x"0E",x"BE",
x"20",x"17",x"7B",x"81",x"FE",x"31",x"20",x"04",x"35",x"37",x"18",x"0E",x"D5",x"C5",
x"CD",x"CB",x"D2",x"F1",x"D1",x"47",x"79",x"3D",x"CD",x"9F",x"D3",x"B7",x"08",x"B7",
x"0D",x"1D",x"D5",x"C5",x"E5",x"F5",x"28",x"02",x"06",x"01",x"C5",x"CD",x"92",x"D5",
x"C1",x"11",x"6B",x"0E",x"1A",x"67",x"69",x"CD",x"87",x"D3",x"E5",x"08",x"30",x"02",
x"2B",x"04",x"1A",x"90",x"4F",x"06",x"00",x"54",x"5D",x"2B",x"28",x"02",x"ED",x"B8",
x"E1",x"01",x"C0",x"FF",x"09",x"46",x"F1",x"20",x"02",x"06",x"20",x"78",x"12",x"E1",
x"C1",x"D1",x"2B",x"20",x"C1",x"ED",x"43",x"49",x"0E",x"C9",x"05",x"20",x"08",x"0D",
x"C8",x"79",x"CD",x"9F",x"D3",x"D0",x"47",x"ED",x"43",x"49",x"0E",x"CD",x"9C",x"D3",
x"B8",x"D8",x"08",x"7E",x"E6",x"7F",x"90",x"38",x"30",x"E5",x"F5",x"D5",x"C5",x"CD",
x"42",x"D5",x"C1",x"D1",x"60",x"69",x"CD",x"87",x"D3",x"08",x"7E",x"30",x"01",x"12",
x"54",x"5D",x"23",x"F1",x"C5",x"28",x"05",x"4F",x"06",x"00",x"ED",x"B0",x"3E",x"20",
x"12",x"C1",x"0C",x"06",x"01",x"E1",x"CB",x"7E",x"23",x"37",x"20",x"CC",x"2B",x"35",
x"C9",x"2B",x"35",x"CB",x"BE",x"79",x"C3",x"1E",x"D3",x"CB",x"FE",x"79",x"FE",x"19",
x"28",x"3F",x"23",x"7E",x"B7",x"C8",x"C5",x"CD",x"09",x"D5",x"C1",x"C5",x"3E",x"19",
x"91",x"21",x"66",x"0E",x"11",x"67",x"0E",x"D5",x"06",x"00",x"4F",x"ED",x"B8",x"13",
x"EB",x"71",x"E1",x"CB",x"BE",x"1F",x"CB",x"19",x"1F",x"CB",x"19",x"47",x"21",x"BF",
x"06",x"11",x"FF",x"06",x"ED",x"B8",x"06",x"40",x"3E",x"20",x"13",x"12",x"10",x"FC",
x"C1",x"21",x"4E",x"0E",x"7E",x"91",x"D8",x"34",x"C9",x"3E",x"01",x"CD",x"1E",x"D3",
x"01",x"18",x"01",x"ED",x"43",x"49",x"0E",x"C9",x"F5",x"4F",x"21",x"4E",x"0E",x"96",
x"CC",x"39",x"D0",x"30",x"01",x"35",x"CD",x"E0",x"D4",x"C1",x"78",x"CD",x"9F",x"D3",
x"E5",x"68",x"26",x"01",x"CD",x"87",x"D3",x"EB",x"21",x"40",x"00",x"19",x"3E",x"18",
x"90",x"F5",x"28",x"0B",x"0E",x"00",x"1F",x"CB",x"19",x"1F",x"CB",x"19",x"47",x"ED",
x"B0",x"06",x"40",x"2B",x"36",x"20",x"10",x"FB",x"F1",x"4F",x"E1",x"54",x"5D",x"23",
x"28",x"02",x"ED",x"B0",x"AF",x"12",x"C9",x"79",x"FE",x"18",x"28",x"A9",x"0C",x"06",
x"01",x"ED",x"43",x"49",x"0E",x"C9",x"ED",x"4B",x"49",x"0E",x"B7",x"0D",x"79",x"C4",
x"9F",x"D3",x"38",x"F8",x"0C",x"06",x"01",x"ED",x"43",x"49",x"0E",x"C9",x"2A",x"49",
x"0E",x"25",x"2D",x"7C",x"87",x"87",x"65",x"CB",x"1C",x"1F",x"CB",x"1C",x"1F",x"6F",
x"7C",x"C6",x"01",x"67",x"22",x"4B",x"0E",x"C9",x"3A",x"49",x"0E",x"C6",x"4F",x"6F",
x"3E",x"0E",x"CE",x"00",x"67",x"7E",x"07",x"B7",x"CB",x"1F",x"C9",x"11",x"40",x"00",
x"D9",x"7E",x"D9",x"A1",x"A8",x"77",x"19",x"D9",x"23",x"10",x"F6",x"C9",x"D9",x"7E",
x"D9",x"57",x"0F",x"0F",x"0F",x"0F",x"AA",x"A1",x"5F",x"E6",x"0F",x"AA",x"A1",x"A8",
x"77",x"2C",x"AB",x"77",x"11",x"3F",x"00",x"19",x"D9",x"23",x"10",x"E5",x"C9",x"D9",
x"7E",x"D9",x"17",x"5F",x"9F",x"57",x"CB",x"13",x"9F",x"AA",x"E6",x"55",x"AA",x"A1",
x"A8",x"77",x"2C",x"CB",x"13",x"9F",x"57",x"CB",x"13",x"9F",x"AA",x"E6",x"55",x"AA",
x"A1",x"A8",x"77",x"2C",x"CB",x"13",x"9F",x"57",x"CB",x"13",x"9F",x"AA",x"E6",x"55",
x"AA",x"A1",x"A8",x"77",x"2C",x"CB",x"13",x"9F",x"57",x"CB",x"13",x"9F",x"AA",x"E6",
x"55",x"AA",x"A1",x"A8",x"77",x"11",x"3D",x"00",x"19",x"D9",x"23",x"10",x"BB",x"C9",
x"08",x"CD",x"59",x"D4",x"E5",x"08",x"4F",x"06",x"00",x"69",x"60",x"29",x"29",x"09",
x"29",x"CB",x"79",x"01",x"74",x"C4",x"28",x"03",x"01",x"40",x"02",x"09",x"06",x"0A",
x"D9",x"3A",x"96",x"0E",x"47",x"3A",x"95",x"0E",x"4F",x"E1",x"C3",x"68",x"0E",x"08",
x"CD",x"05",x"CC",x"32",x"96",x"0E",x"CD",x"0D",x"CC",x"A8",x"32",x"95",x"0E",x"08",
x"C9",x"05",x"3A",x"73",x"0B",x"B7",x"28",x"05",x"CB",x"20",x"3D",x"20",x"FB",x"0D",
x"79",x"87",x"87",x"81",x"87",x"67",x"AF",x"CB",x"3C",x"1F",x"37",x"CB",x"1C",x"1F",
x"B0",x"6F",x"C9",x"CD",x"59",x"D4",x"11",x"6D",x"0E",x"3A",x"6C",x"0E",x"4F",x"06",
x"0A",x"C5",x"E5",x"06",x"00",x"ED",x"B0",x"E1",x"0E",x"40",x"09",x"C1",x"10",x"F3",
x"C9",x"CD",x"59",x"D4",x"11",x"6D",x"0E",x"3A",x"6C",x"0E",x"4F",x"06",x"0A",x"EB",
x"C5",x"D5",x"06",x"00",x"ED",x"B0",x"EB",x"E1",x"0E",x"40",x"09",x"C1",x"10",x"F1",
x"C9",x"CD",x"59",x"D4",x"3A",x"96",x"0E",x"08",x"3E",x"3F",x"95",x"E6",x"3F",x"28",
x"18",x"4F",x"7D",x"06",x"0A",x"E6",x"3F",x"B5",x"6F",x"08",x"77",x"54",x"5D",x"1C",
x"C5",x"06",x"00",x"ED",x"B0",x"C1",x"EB",x"08",x"10",x"ED",x"C9",x"11",x"40",x"00",
x"06",x"0A",x"3A",x"96",x"0E",x"77",x"19",x"10",x"FC",x"C9",x"79",x"FE",x"18",x"28",
x"14",x"06",x"01",x"CD",x"59",x"D4",x"EB",x"21",x"80",x"B9",x"B7",x"ED",x"52",x"44",
x"4D",x"21",x"80",x"02",x"19",x"ED",x"B0",x"21",x"80",x"B9",x"11",x"81",x"B9",x"01",
x"7F",x"02",x"3A",x"96",x"0E",x"77",x"ED",x"B0",x"C9",x"3E",x"18",x"91",x"28",x"EB",
x"4F",x"87",x"87",x"81",x"87",x"47",x"AF",x"CB",x"38",x"1F",x"CB",x"38",x"1F",x"4F",
x"21",x"7F",x"B9",x"11",x"FF",x"BB",x"ED",x"B8",x"23",x"54",x"5D",x"13",x"18",x"D5",
x"3A",x"6C",x"0E",x"4F",x"06",x"0A",x"C5",x"E5",x"D5",x"06",x"00",x"ED",x"B0",x"0E",
x"40",x"E1",x"09",x"EB",x"E1",x"09",x"C1",x"10",x"EF",x"C9",x"28",x"1E",x"E5",x"C5",
x"5F",x"3A",x"73",x"0B",x"B7",x"28",x"05",x"CB",x"23",x"3D",x"20",x"FB",x"CD",x"59",
x"D4",x"4B",x"54",x"3A",x"6C",x"0E",x"85",x"5F",x"EB",x"CD",x"2E",x"D5",x"C1",x"E1",
x"46",x"CB",x"78",x"28",x"11",x"C5",x"CB",x"B8",x"CD",x"59",x"D4",x"EB",x"C1",x"0C",
x"06",x"01",x"CD",x"59",x"D4",x"C3",x"2A",x"D5",x"CD",x"59",x"D4",x"0E",x"0A",x"11",
x"40",x"00",x"3A",x"6C",x"0E",x"47",x"3A",x"96",x"0E",x"E5",x"77",x"23",x"10",x"FC",
x"E1",x"19",x"0D",x"20",x"EF",x"C9",x"F5",x"7E",x"E6",x"7F",x"90",x"28",x"35",x"5F",
x"3A",x"73",x"0B",x"B7",x"28",x"05",x"CB",x"23",x"3D",x"20",x"FB",x"E5",x"C5",x"46",
x"CB",x"B8",x"CD",x"59",x"D4",x"2B",x"4B",x"06",x"00",x"EB",x"3A",x"6C",x"0E",x"6F",
x"60",x"19",x"EB",x"06",x"0A",x"C5",x"E5",x"D5",x"06",x"00",x"ED",x"B8",x"0E",x"40",
x"E1",x"09",x"EB",x"E1",x"09",x"C1",x"10",x"EF",x"C1",x"E1",x"F1",x"28",x"A7",x"EB",
x"C5",x"CD",x"59",x"D4",x"C1",x"EB",x"0D",x"2B",x"46",x"CB",x"B8",x"CD",x"59",x"D4",
x"C3",x"2A",x"D5",x"04",x"2D",x"D6",x"18",x"D6",x"2C",x"D6",x"12",x"D6",x"3E",x"1E",
x"32",x"65",x"0B",x"3E",x"03",x"32",x"67",x"0B",x"AF",x"32",x"66",x"0B",x"21",x"51",
x"0B",x"11",x"52",x"0B",x"01",x"13",x"00",x"77",x"ED",x"B0",x"21",x"E5",x"0B",x"11",
x"E6",x"0B",x"0E",x"09",x"77",x"ED",x"B0",x"C9",x"3A",x"E5",x"0B",x"4F",x"AF",x"C9",
x"21",x"E5",x"0B",x"7E",x"B7",x"28",x"FC",x"3A",x"E9",x"0B",x"4F",x"36",x"00",x"3A",
x"16",x"0B",x"B7",x"C8",x"3E",x"F5",x"C9",x"3A",x"66",x"0B",x"E6",x"0B",x"47",x"ED",
x"44",x"A0",x"32",x"66",x"0B",x"CD",x"A5",x"D7",x"21",x"E7",x"0B",x"FD",x"CB",x"06",
x"6E",x"28",x"0D",x"7E",x"B7",x"C0",x"35",x"3E",x"01",x"CD",x"90",x"D7",x"32",x"66",
x"0B",x"C0",x"70",x"3E",x"04",x"CD",x"90",x"D7",x"32",x"E8",x"0B",x"AF",x"CD",x"C7",
x"D6",x"1C",x"28",x"10",x"79",x"32",x"E9",x"0B",x"3E",x"FF",x"32",x"E5",x"0B",x"3A",
x"65",x"0B",x"32",x"EA",x"0B",x"C9",x"7E",x"B7",x"20",x"E6",x"21",x"EA",x"0B",x"CD",
x"C0",x"D6",x"23",x"D4",x"C0",x"D6",x"D0",x"3A",x"EE",x"0B",x"4F",x"ED",x"5B",x"EC",
x"0B",x"21",x"64",x"0B",x"ED",x"52",x"EB",x"28",x"0A",x"B7",x"EB",x"21",x"64",x"0B",
x"ED",x"52",x"EB",x"20",x"09",x"16",x"66",x"A2",x"28",x"04",x"AA",x"A6",x"20",x"11",
x"79",x"A6",x"20",x"0D",x"21",x"5B",x"0B",x"06",x"0A",x"77",x"23",x"10",x"FC",x"32",
x"EB",x"0B",x"C9",x"2F",x"A6",x"77",x"3A",x"67",x"0B",x"32",x"EB",x"0B",x"18",x"9B",
x"7E",x"B7",x"C8",x"35",x"C0",x"37",x"C9",x"C4",x"A5",x"D7",x"FD",x"CB",x"06",x"9E",
x"FD",x"CB",x"07",x"A6",x"FD",x"CB",x"07",x"86",x"FD",x"CB",x"06",x"AE",x"21",x"E6",
x"0B",x"11",x"0A",x"00",x"D9",x"21",x"65",x"0B",x"11",x"5B",x"0B",x"1B",x"2B",x"D9",
x"1D",x"F8",x"D9",x"1A",x"47",x"AE",x"2F",x"A6",x"77",x"A8",x"28",x"F1",x"47",x"ED",
x"44",x"A0",x"47",x"AE",x"77",x"78",x"22",x"EC",x"0B",x"32",x"EE",x"0B",x"3E",x"50",
x"D6",x"0A",x"CB",x"38",x"30",x"FA",x"D9",x"83",x"5F",x"3A",x"E8",x"0B",x"47",x"3A",
x"66",x"0B",x"A8",x"47",x"E5",x"CD",x"47",x"D7",x"E1",x"3A",x"68",x"0B",x"3C",x"C8",
x"7E",x"B7",x"79",x"28",x"15",x"3A",x"11",x"0B",x"E6",x"F0",x"F6",x"07",x"D3",x"03",
x"DB",x"58",x"E6",x"18",x"28",x"0A",x"AF",x"32",x"16",x"0B",x"18",x"04",x"FE",x"10",
x"28",x"03",x"36",x"00",x"C9",x"35",x"1E",x"FF",x"C9",x"21",x"84",x"D7",x"E5",x"21",
x"5F",x"D8",x"CB",x"50",x"C0",x"CB",x"40",x"28",x"1F",x"21",x"BF",x"D7",x"19",x"7E",
x"FE",x"61",x"38",x"16",x"FE",x"7B",x"38",x"08",x"FE",x"90",x"38",x"0E",x"FE",x"99",
x"30",x"0A",x"21",x"0F",x"D8",x"CB",x"48",x"C8",x"21",x"BF",x"D7",x"C9",x"21",x"0F",
x"D8",x"CB",x"48",x"C0",x"21",x"AF",x"D8",x"CB",x"58",x"C0",x"E1",x"21",x"BF",x"D7",
x"19",x"4E",x"79",x"FE",x"FF",x"C0",x"32",x"16",x"0B",x"0E",x"1B",x"C9",x"FD",x"CB",
x"07",x"66",x"C0",x"3E",x"02",x"FD",x"CB",x"06",x"5E",x"C0",x"FD",x"CB",x"07",x"46",
x"3E",x"08",x"C0",x"AF",x"C9",x"3A",x"11",x"0B",x"E6",x"F0",x"4F",x"21",x"51",x"0B",
x"E5",x"FD",x"E1",x"06",x"0A",x"79",x"D3",x"03",x"DB",x"58",x"2F",x"77",x"0C",x"23",
x"10",x"F5",x"C9",x"34",x"37",x"72",x"75",x"66",x"6A",x"76",x"6D",x"2A",x"2A",x"31",
x"94",x"71",x"70",x"61",x"91",x"79",x"2D",x"13",x"F3",x"92",x"93",x"40",x"96",x"3C",
x"98",x"2A",x"20",x"04",x"E4",x"36",x"2A",x"7A",x"5B",x"68",x"0D",x"6E",x"2A",x"01",
x"E1",x"30",x"97",x"3B",x"95",x"5C",x"90",x"2A",x"1B",x"06",x"E6",x"32",x"39",x"77",
x"6F",x"73",x"6C",x"78",x"2E",x"18",x"F8",x"33",x"38",x"65",x"69",x"64",x"6B",x"63",
x"2C",x"05",x"E5",x"35",x"5E",x"74",x"5D",x"67",x"08",x"62",x"2A",x"16",x"43",x"21",
x"3D",x"52",x"55",x"46",x"4A",x"56",x"4D",x"2A",x"2A",x"27",x"84",x"51",x"50",x"41",
x"81",x"59",x"5F",x"13",x"F3",x"82",x"83",x"60",x"86",x"3E",x"88",x"2A",x"20",x"04",
x"E4",x"2F",x"23",x"5A",x"7B",x"48",x"0D",x"4E",x"2A",x"01",x"E1",x"26",x"87",x"24",
x"85",x"7C",x"80",x"2A",x"1B",x"06",x"E6",x"22",x"29",x"57",x"4F",x"53",x"4C",x"58",
x"3A",x"18",x"F8",x"2B",x"28",x"45",x"49",x"44",x"4B",x"43",x"3F",x"05",x"E5",x"25",
x"7E",x"54",x"7D",x"47",x"07",x"42",x"2A",x"16",x"49",x"8B",x"9C",x"12",x"15",x"06",
x"0A",x"16",x"0D",x"2A",x"2A",x"99",x"DC",x"11",x"10",x"01",x"D9",x"19",x"1F",x"13",
x"F3",x"DA",x"DB",x"00",x"DE",x"3C",x"98",x"2A",x"20",x"04",x"E4",x"8C",x"8E",x"1A",
x"1B",x"08",x"0D",x"0E",x"2A",x"01",x"E1",x"89",x"DF",x"3B",x"DD",x"1C",x"CF",x"2A",
x"FF",x"06",x"E6",x"8A",x"9D",x"17",x"0F",x"13",x"0C",x"18",x"2E",x"18",x"F8",x"9A",
x"8D",x"05",x"09",x"04",x"0B",x"03",x"2C",x"05",x"E5",x"9B",x"1E",x"14",x"1D",x"07",
x"08",x"02",x"2A",x"16",x"53",x"A4",x"A7",x"C2",x"C5",x"B6",x"BA",x"C6",x"BD",x"2A",
x"2A",x"A1",x"D4",x"C1",x"C0",x"B1",x"D1",x"C9",x"AD",x"13",x"F3",x"D2",x"D3",x"B0",
x"D6",x"AC",x"D8",x"2A",x"20",x"04",x"E4",x"A6",x"AA",x"CA",x"CB",x"B8",x"0D",x"BE",
x"2A",x"01",x"E1",x"A0",x"D7",x"AB",x"D5",x"CC",x"D0",x"2A",x"1B",x"06",x"E6",x"A2",
x"A9",x"C7",x"BF",x"C3",x"BC",x"C8",x"AE",x"18",x"F8",x"A3",x"A8",x"B5",x"B9",x"B4",
x"BB",x"B3",x"AF",x"05",x"E5",x"A5",x"CE",x"C4",x"CD",x"B7",x"08",x"B2",x"2A",x"16",
x"4C",x"03",x"29",x"D9",x"0C",x"D9",x"06",x"D9",x"21",x"0C",x"D9",x"C3",x"6D",x"C5",
x"3A",x"16",x"0B",x"3C",x"3E",x"F5",x"C8",x"DB",x"59",x"07",x"30",x"F4",x"F3",x"79",
x"D3",x"01",x"3A",x"13",x"0B",x"E6",x"7F",x"D3",x"06",x"F6",x"80",x"D3",x"06",x"FB",
x"AF",x"C9",x"04",x"33",x"D9",x"60",x"D9",x"60",x"D9",x"61",x"D9",x"3A",x"14",x"0B",
x"3C",x"C0",x"3A",x"16",x"0B",x"3C",x"28",x"08",x"3A",x"EF",x"0B",x"3D",x"32",x"EF",
x"0B",x"C0",x"32",x"14",x"0B",x"32",x"EF",x"0B",x"3A",x"10",x"0B",x"F6",x"08",x"32",
x"10",x"0B",x"3A",x"12",x"0B",x"E6",x"CF",x"32",x"12",x"0B",x"D3",x"05",x"3E",x"F5",
x"C9",x"3A",x"15",x"0B",x"3C",x"28",x"07",x"3A",x"EF",x"0B",x"D6",x"02",x"30",x"F3",
x"AF",x"32",x"14",x"0B",x"3A",x"16",x"0B",x"3C",x"28",x"CE",x"78",x"B7",x"20",x"05",
x"CD",x"46",x"D9",x"AF",x"C9",x"32",x"EF",x"0B",x"79",x"E6",x"0F",x"07",x"07",x"4F",
x"3A",x"13",x"0B",x"E6",x"C3",x"B1",x"32",x"13",x"0B",x"D3",x"06",x"7A",x"E6",x"0F",
x"F6",x"10",x"57",x"3A",x"12",x"0B",x"E6",x"C0",x"B2",x"32",x"12",x"0B",x"D3",x"05",
x"7B",x"D3",x"04",x"3E",x"FF",x"32",x"14",x"0B",x"32",x"71",x"0B",x"3A",x"10",x"0B",
x"E6",x"F7",x"32",x"10",x"0B",x"AF",x"C9",x"06",x"E7",x"D9",x"D2",x"D9",x"D7",x"D9",
x"C8",x"D9",x"CD",x"D9",x"DC",x"D9",x"21",x"E2",x"F3",x"18",x"12",x"21",x"E7",x"F3",
x"18",x"0D",x"21",x"D8",x"F3",x"18",x"08",x"21",x"DD",x"F3",x"18",x"03",x"21",x"EC",
x"F3",x"C3",x"F0",x"FF",x"21",x"F1",x"F3",x"18",x"F8",x"C9",x"28",x"63",x"29",x"20",
x"49",x"53",x"4C",x"21",x"00",x"17",x"E5",x"DD",x"E1",x"3A",x"21",x"0B",x"B7",x"C2",
x"D3",x"DA",x"01",x"EF",x"02",x"77",x"ED",x"A1",x"EA",x"FF",x"D9",x"22",x"20",x"17",
x"22",x"22",x"17",x"21",x"5B",x"FB",x"11",x"08",x"00",x"01",x"27",x"00",x"ED",x"B0",
x"CD",x"10",x"DE",x"11",x"15",x"DC",x"F7",x"0C",x"3E",x"02",x"32",x"4F",x"0B",x"DD",
x"36",x"05",x"00",x"01",x"03",x"03",x"3E",x"0C",x"C5",x"F5",x"F7",x"03",x"CD",x"F2",
x"DB",x"F1",x"F5",x"CD",x"0C",x"DC",x"CD",x"F2",x"DB",x"CD",x"93",x"FE",x"F1",x"C1",
x"04",x"0C",x"0C",x"D6",x"02",x"30",x"E5",x"01",x"15",x"0D",x"F7",x"03",x"CD",x"F2",
x"DB",x"01",x"12",x"0B",x"F7",x"03",x"21",x"FF",x"DB",x"46",x"23",x"7E",x"CD",x"9A",
x"FE",x"E5",x"C5",x"CD",x"D8",x"E6",x"E6",x"03",x"28",x"F9",x"C1",x"E1",x"32",x"4D",
x"0B",x"0D",x"20",x"FD",x"10",x"E8",x"F7",x"93",x"0C",x"20",x"DA",x"F7",x"91",x"0E",
x"01",x"F7",x"04",x"32",x"4F",x"0B",x"CD",x"18",x"FC",x"CD",x"79",x"FE",x"32",x"54",
x"56",x"20",x"43",x"4F",x"4D",x"50",x"55",x"54",x"45",x"52",x"20",x"42",x"41",x"53",
x"49",x"43",x"20",x"31",x"2E",x"32",x"0D",x"0A",x"43",x"6F",x"70",x"79",x"72",x"69",
x"67",x"68",x"74",x"20",x"31",x"39",x"38",x"35",x"20",x"56",x"49",x"44",x"45",x"4F",
x"54",x"4F",x"4E",x"0D",x"0A",x"0D",x"0A",x"CD",x"4C",x"EC",x"CD",x"C1",x"FE",x"CD",
x"1B",x"FA",x"CD",x"79",x"FE",x"0F",x"20",x"62",x"79",x"74",x"65",x"73",x"20",x"66",
x"72",x"65",x"65",x"0D",x"0A",x"0D",x"0A",x"AF",x"32",x"21",x"0B",x"CD",x"FC",x"DC",
x"31",x"AC",x"16",x"21",x"03",x"17",x"7E",x"B7",x"36",x"00",x"C4",x"10",x"DE",x"DD",
x"36",x"05",x"20",x"DD",x"CB",x"00",x"96",x"DD",x"CB",x"00",x"4E",x"20",x"0A",x"CD",
x"18",x"FC",x"CD",x"79",x"FE",x"03",x"6F",x"6B",x"0B",x"DD",x"CB",x"00",x"8E",x"CD",
x"93",x"FE",x"CD",x"4F",x"FF",x"FE",x"F5",x"CA",x"A3",x"FF",x"FE",x"EC",x"28",x"E3",
x"CD",x"19",x"DC",x"5D",x"54",x"23",x"CD",x"14",x"F9",x"38",x"0D",x"7E",x"FE",x"A8",
x"28",x"03",x"3C",x"20",x"3C",x"CD",x"1B",x"FA",x"18",x"DC",x"17",x"38",x"34",x"46",
x"FD",x"7E",x"08",x"FE",x"40",x"38",x"2C",x"FE",x"44",x"30",x"28",x"FD",x"7E",x"06",
x"B7",x"28",x"22",x"7E",x"23",x"FE",x"20",x"28",x"FA",x"2B",x"EB",x"7E",x"23",x"C6",
x"02",x"ED",x"52",x"85",x"4F",x"CD",x"C3",x"FA",x"EB",x"2B",x"72",x"2B",x"73",x"2B",
x"71",x"22",x"0C",x"17",x"CD",x"AF",x"DC",x"18",x"A5",x"EB",x"CD",x"1B",x"FA",x"4E",
x"AF",x"77",x"2B",x"77",x"2B",x"0C",x"0C",x"71",x"22",x"0C",x"17",x"23",x"DD",x"CB",
x"00",x"46",x"C4",x"4D",x"DE",x"DD",x"CB",x"02",x"86",x"23",x"23",x"D9",x"D9",x"CD",
x"9D",x"FF",x"FD",x"22",x"1A",x"17",x"7E",x"FE",x"FE",x"30",x"2E",x"23",x"FE",x"20",
x"28",x"F6",x"FE",x"CA",x"DA",x"BC",x"E3",x"F5",x"D9",x"2F",x"87",x"C6",x"67",x"6F",
x"26",x"C0",x"7E",x"2C",x"66",x"6F",x"F1",x"FE",x"FB",x"DC",x"43",x"FC",x"31",x"AC",
x"16",x"E9",x"CD",x"43",x"FC",x"D9",x"78",x"D9",x"FE",x"FD",x"28",x"C8",x"DA",x"5A",
x"FD",x"2A",x"0C",x"17",x"4E",x"AF",x"47",x"09",x"B6",x"20",x"A9",x"FD",x"7E",x"00",
x"FE",x"2B",x"28",x"0E",x"FE",x"06",x"28",x"0A",x"DD",x"CB",x"00",x"56",x"CA",x"DA",
x"DA",x"C3",x"0E",x"E1",x"FD",x"5E",x"03",x"FD",x"56",x"04",x"21",x"31",x"18",x"ED",
x"52",x"38",x"E9",x"4F",x"06",x"00",x"FD",x"09",x"FD",x"22",x"1A",x"17",x"18",x"D3",
x"CD",x"79",x"FE",x"08",x"56",x"49",x"44",x"45",x"4F",x"54",x"4F",x"4E",x"C9",x"0C",
x"54",x"56",x"20",x"20",x"43",x"4F",x"4D",x"50",x"55",x"54",x"45",x"52",x"3D",x"F8",
x"F5",x"CD",x"C7",x"FE",x"F1",x"18",x"F7",x"01",x"44",x"54",x"51",x"FD",x"E5",x"EB",
x"FD",x"21",x"35",x"17",x"01",x"00",x"00",x"13",x"21",x"6E",x"DE",x"3E",x"FE",x"08",
x"FD",x"23",x"ED",x"53",x"1C",x"17",x"CD",x"BF",x"FB",x"FD",x"77",x"00",x"3C",x"28",
x"66",x"78",x"B7",x"28",x"04",x"FE",x"3A",x"20",x"0A",x"1A",x"FE",x"22",x"20",x"05",
x"48",x"47",x"13",x"18",x"DF",x"CD",x"BF",x"FB",x"13",x"B7",x"28",x"0E",x"B8",x"20",
x"0B",x"41",x"0E",x"00",x"FE",x"22",x"28",x"C8",x"3E",x"FD",x"18",x"28",x"04",x"05",
x"20",x"C6",x"AE",x"87",x"20",x"25",x"23",x"30",x"E0",x"08",x"48",x"FE",x"A6",x"28",
x"08",x"FE",x"A5",x"28",x"04",x"FE",x"A3",x"20",x"02",x"D6",x"08",x"FE",x"FD",x"28",
x"09",x"FE",x"FB",x"38",x"05",x"47",x"20",x"02",x"06",x"3A",x"FD",x"77",x"00",x"18",
x"97",x"ED",x"5B",x"1C",x"17",x"CB",x"7E",x"23",x"28",x"FB",x"08",x"3D",x"08",x"7E",
x"3C",x"28",x"86",x"18",x"AC",x"FD",x"E5",x"E1",x"23",x"77",x"11",x"35",x"17",x"B7",
x"ED",x"52",x"EB",x"73",x"FD",x"E1",x"C9",x"22",x"1C",x"17",x"C5",x"CD",x"45",x"DD",
x"D4",x"E6",x"DC",x"C1",x"04",x"C8",x"06",x"00",x"CD",x"C9",x"DC",x"EB",x"2A",x"1C",
x"17",x"ED",x"B0",x"18",x"33",x"CD",x"FC",x"DC",x"CD",x"8E",x"FC",x"C5",x"E5",x"CD",
x"41",x"DD",x"D1",x"E5",x"B7",x"ED",x"52",x"4D",x"44",x"D1",x"E1",x"E5",x"19",x"EB",
x"03",x"ED",x"B8",x"23",x"C1",x"C9",x"4E",x"06",x"00",x"E5",x"09",x"E5",x"CD",x"41",
x"DD",x"D1",x"B7",x"ED",x"52",x"4D",x"44",x"EB",x"D1",x"D5",x"03",x"ED",x"B0",x"E1",
x"E5",x"D5",x"C5",x"FD",x"2A",x"19",x"0B",x"21",x"00",x"00",x"FD",x"75",x"00",x"22",
x"0E",x"17",x"22",x"14",x"17",x"21",x"94",x"F0",x"22",x"24",x"17",x"21",x"09",x"17",
x"75",x"22",x"0A",x"17",x"2A",x"22",x"17",x"22",x"12",x"17",x"CD",x"41",x"DD",x"23",
x"22",x"26",x"17",x"C1",x"D1",x"E1",x"C9",x"F5",x"23",x"5E",x"23",x"56",x"23",x"E5",
x"EB",x"CD",x"19",x"FF",x"E1",x"CD",x"DD",x"FE",x"F1",x"D0",x"C3",x"8E",x"FE",x"21",
x"FF",x"FF",x"EB",x"2A",x"22",x"17",x"01",x"00",x"00",x"09",x"4E",x"0C",x"0D",x"37",
x"C8",x"D5",x"23",x"5E",x"23",x"56",x"2B",x"2B",x"E3",x"B7",x"ED",x"52",x"19",x"EB",
x"E1",x"C8",x"30",x"E9",x"C9",x"CF",x"0A",x"DD",x"CB",x"00",x"56",x"C2",x"B1",x"DB",
x"DD",x"CB",x"00",x"D6",x"2A",x"0E",x"17",x"7C",x"B5",x"28",x"EC",x"22",x"0C",x"17",
x"2A",x"10",x"17",x"C3",x"81",x"DB",x"0E",x"40",x"B1",x"18",x"03",x"0E",x"20",x"AF",
x"F5",x"CD",x"EE",x"FB",x"F1",x"20",x"05",x"79",x"FE",x"20",x"16",x"F6",x"37",x"08",
x"D9",x"78",x"D9",x"21",x"00",x"00",x"11",x"FF",x"FF",x"FE",x"FD",x"30",x"2E",x"18",
x"11",x"D9",x"78",x"D9",x"FE",x"A4",x"28",x"07",x"08",x"DA",x"B1",x"DB",x"C3",x"DA",
x"DA",x"CD",x"43",x"FC",x"CD",x"FB",x"DD",x"14",x"20",x"08",x"FE",x"A2",x"C2",x"5A",
x"FD",x"11",x"00",x"01",x"15",x"D5",x"FE",x"A2",x"20",x"06",x"CD",x"43",x"FC",x"CD",
x"FB",x"DD",x"E1",x"D5",x"CD",x"44",x"DD",x"D1",x"7E",x"B7",x"28",x"CB",x"23",x"4E",
x"23",x"46",x"2B",x"2B",x"EB",x"ED",x"42",x"09",x"EB",x"38",x"BE",x"D5",x"08",x"30",
x"05",x"CD",x"2D",x"DD",x"18",x"04",x"CD",x"E6",x"DC",x"B7",x"08",x"CD",x"9D",x"FF",
x"D1",x"18",x"DB",x"11",x"FF",x"FF",x"FE",x"02",x"C0",x"CD",x"C3",x"FA",x"EB",x"C3",
x"43",x"FC",x"21",x"DA",x"DA",x"E5",x"DD",x"CB",x"00",x"86",x"2A",x"20",x"17",x"22",
x"22",x"17",x"36",x"00",x"C3",x"FC",x"DC",x"2A",x"22",x"17",x"FE",x"02",x"CC",x"DE",
x"FB",x"CD",x"FC",x"DC",x"CD",x"3E",x"FC",x"DD",x"CB",x"00",x"D6",x"AF",x"C3",x"C2",
x"DB",x"CD",x"EC",x"FB",x"DD",x"71",x"06",x"FE",x"E3",x"28",x"0B",x"FE",x"C1",x"C2",
x"5A",x"FD",x"DD",x"CB",x"00",x"86",x"18",x"04",x"DD",x"CB",x"00",x"C6",x"C3",x"AE",
x"DB",x"DD",x"CB",x"00",x"56",x"C8",x"3A",x"06",x"17",x"32",x"05",x"17",x"E5",x"5E",
x"23",x"56",x"EB",x"3E",x"3C",x"CD",x"9A",x"FE",x"06",x"00",x"CD",x"1B",x"FF",x"E1",
x"3E",x"3E",x"C3",x"9A",x"FE",x"FF",x"A1",x"BA",x"52",x"45",x"CD",x"44",x"41",x"54",
x"C1",x"43",x"4C",x"4F",x"53",x"C5",x"43",x"4C",x"D3",x"43",x"4F",x"4E",x"54",x"49",
x"4E",x"55",x"C5",x"44",x"45",x"C6",x"44",x"45",x"4C",x"45",x"54",x"C5",x"44",x"49",
x"CD",x"45",x"4C",x"53",x"C5",x"45",x"4E",x"C4",x"46",x"4F",x"D2",x"47",x"45",x"D4",
x"47",x"4F",x"53",x"55",x"C2",x"47",x"4F",x"54",x"CF",x"47",x"52",x"41",x"50",x"48",
x"49",x"43",x"D3",x"49",x"C6",x"49",x"4E",x"50",x"55",x"D4",x"4C",x"45",x"D4",x"4C",
x"49",x"53",x"D4",x"4C",x"4C",x"49",x"53",x"D4",x"4C",x"4F",x"41",x"C4",x"4C",x"4F",
x"4D",x"45",x"CD",x"4E",x"45",x"D7",x"4E",x"45",x"58",x"D4",x"4F",x"CB",x"4F",x"CE",
x"4F",x"50",x"45",x"CE",x"4F",x"55",x"54",x"50",x"55",x"D4",x"4F",x"55",x"D4",x"50",
x"4C",x"4F",x"D4",x"50",x"4F",x"4B",x"C5",x"50",x"52",x"49",x"4E",x"D4",x"52",x"41",
x"4E",x"44",x"4F",x"4D",x"49",x"5A",x"C5",x"52",x"45",x"41",x"C4",x"52",x"45",x"53",
x"54",x"4F",x"52",x"C5",x"52",x"45",x"54",x"55",x"52",x"CE",x"52",x"55",x"CE",x"53",
x"41",x"56",x"C5",x"53",x"45",x"D4",x"53",x"4F",x"55",x"4E",x"C4",x"53",x"54",x"4F",
x"D0",x"54",x"52",x"41",x"43",x"C5",x"56",x"45",x"52",x"49",x"46",x"D9",x"45",x"58",
x"D4",x"4C",x"50",x"52",x"49",x"4E",x"D4",x"A1",x"A1",x"A1",x"A1",x"A1",x"A1",x"41",
x"4E",x"C4",x"43",x"48",x"41",x"52",x"41",x"43",x"54",x"45",x"D2",x"44",x"45",x"4C",
x"41",x"D9",x"44",x"55",x"52",x"41",x"54",x"49",x"4F",x"CE",x"49",x"4E",x"4B",x"45",
x"59",x"A4",x"49",x"4E",x"CB",x"4D",x"4F",x"44",x"C5",x"4E",x"4F",x"D4",x"4F",x"46",
x"C6",x"4F",x"52",x"C4",x"4F",x"D2",x"50",x"41",x"49",x"4E",x"D4",x"50",x"41",x"4C",
x"45",x"54",x"54",x"C5",x"50",x"41",x"50",x"45",x"D2",x"50",x"49",x"54",x"43",x"C8",
x"50",x"52",x"4F",x"4D",x"50",x"D4",x"52",x"41",x"54",x"C5",x"53",x"54",x"45",x"D0",
x"53",x"54",x"59",x"4C",x"C5",x"54",x"41",x"C2",x"54",x"48",x"45",x"CE",x"54",x"CF",
x"56",x"4F",x"4C",x"55",x"4D",x"C5",x"58",x"4F",x"D2",x"41",x"54",x"CE",x"41",x"D4",
x"55",x"53",x"49",x"4E",x"C7",x"42",x"4F",x"52",x"44",x"45",x"D2",x"A1",x"A1",x"A1",
x"A1",x"A1",x"AA",x"A3",x"3D",x"BE",x"3E",x"BC",x"AC",x"3D",x"BC",x"AD",x"AF",x"BB",
x"DE",x"3E",x"BD",x"3C",x"BE",x"BE",x"3C",x"BD",x"BD",x"BC",x"AB",x"A6",x"A8",x"A9",
x"FF",x"20",x"6D",x"69",x"73",x"73",x"69",x"6E",x"E7",x"72",x"67",x"75",x"6D",x"65",
x"6E",x"F4",x"42",x"61",x"64",x"A0",x"4E",x"6F",x"A0",x"43",x"61",x"6E",x"6E",x"6F",
x"74",x"A0",x"D9",x"7E",x"FE",x"FD",x"D2",x"81",x"DB",x"23",x"18",x"F7",x"F7",x"05",
x"D7",x"C3",x"B1",x"DB",x"E6",x"81",x"FE",x"01",x"C2",x"5A",x"FD",x"DD",x"CB",x"00",
x"56",x"28",x"1F",x"D9",x"E5",x"D5",x"D9",x"E1",x"2B",x"CB",x"7E",x"28",x"35",x"CB",
x"BE",x"CB",x"D6",x"23",x"ED",x"5B",x"0C",x"17",x"73",x"23",x"72",x"23",x"D1",x"73",
x"23",x"72",x"23",x"22",x"26",x"17",x"D9",x"0E",x"01",x"0D",x"3E",x"0C",x"7E",x"FE",
x"FE",x"D2",x"4B",x"E0",x"23",x"FE",x"96",x"28",x"F4",x"FE",x"95",x"28",x"EE",x"FE",
x"FD",x"20",x"ED",x"0C",x"0D",x"20",x"E9",x"C3",x"81",x"DB",x"CF",x"0F",x"CD",x"43",
x"FC",x"B7",x"FA",x"5A",x"FD",x"CB",x"47",x"CA",x"5A",x"FD",x"D9",x"79",x"E6",x"88",
x"28",x"EC",x"E6",x"08",x"C4",x"0B",x"F4",x"1B",x"1A",x"EE",x"81",x"32",x"01",x"17",
x"12",x"13",x"3E",x"FF",x"12",x"D5",x"13",x"ED",x"53",x"26",x"17",x"D9",x"CD",x"43",
x"FC",x"DD",x"CB",x"01",x"4E",x"20",x"20",x"FE",x"A8",x"20",x"1C",x"CD",x"16",x"FB",
x"3C",x"28",x"57",x"3D",x"4F",x"E1",x"22",x"26",x"17",x"2B",x"CB",x"86",x"CD",x"C1",
x"F3",x"D9",x"78",x"D9",x"FE",x"A4",x"28",x"B0",x"C3",x"B4",x"DB",x"3E",x"96",x"CD",
x"54",x"FD",x"37",x"D4",x"43",x"FC",x"CD",x"C4",x"FA",x"FA",x"14",x"FB",x"23",x"EB",
x"2A",x"26",x"17",x"73",x"23",x"72",x"23",x"22",x"26",x"17",x"EB",x"CD",x"2B",x"FA",
x"E1",x"34",x"E5",x"C4",x"12",x"F5",x"D9",x"78",x"D9",x"FE",x"A4",x"28",x"DA",x"3E",
x"95",x"CD",x"54",x"FD",x"E1",x"34",x"DD",x"CB",x"01",x"4E",x"20",x"0D",x"FE",x"A8",
x"3E",x"12",x"CC",x"16",x"FB",x"3C",x"CA",x"14",x"FB",x"3D",x"4F",x"C5",x"DF",x"0C",
x"85",x"26",x"CD",x"93",x"F6",x"F2",x"B1",x"FC",x"CD",x"C3",x"FA",x"C1",x"E5",x"CD",
x"BB",x"F3",x"E1",x"2B",x"7D",x"B4",x"20",x"F6",x"18",x"95",x"DD",x"CB",x"02",x"46",
x"CA",x"5A",x"FD",x"C3",x"BB",x"DB",x"21",x"00",x"00",x"22",x"0E",x"17",x"C3",x"DA",
x"DA",x"CD",x"1B",x"FB",x"FE",x"07",x"D2",x"14",x"FB",x"87",x"F5",x"D9",x"78",x"D9",
x"FE",x"A4",x"20",x"16",x"CD",x"BA",x"FA",x"EB",x"FE",x"A4",x"20",x"0E",x"CD",x"BA",
x"FA",x"FE",x"A4",x"20",x"07",x"E5",x"CD",x"BA",x"FA",x"4D",x"44",x"E1",x"E3",x"D5",
x"5C",x"16",x"00",x"21",x"21",x"00",x"19",x"5E",x"23",x"56",x"7A",x"B3",x"CA",x"B1",
x"DB",x"ED",x"53",x"16",x"00",x"D1",x"21",x"B1",x"DB",x"E3",x"EB",x"C3",x"15",x"00",
x"FE",x"03",x"28",x"07",x"E6",x"82",x"C2",x"5A",x"FD",x"CF",x"0E",x"CD",x"2E",x"F4",
x"3E",x"9A",x"CD",x"54",x"FD",x"CD",x"8E",x"FC",x"E5",x"CD",x"A7",x"F0",x"E1",x"E5",
x"CD",x"28",x"FB",x"3E",x"B4",x"CD",x"54",x"FD",x"CD",x"A7",x"F0",x"11",x"EE",x"FF",
x"FD",x"19",x"FE",x"B8",x"28",x"09",x"08",x"21",x"01",x"00",x"CD",x"2B",x"FA",x"08",
x"37",x"D4",x"A4",x"F0",x"FE",x"FD",x"DA",x"5A",x"FD",x"FD",x"E5",x"E1",x"D1",x"2B",
x"72",x"2B",x"73",x"ED",x"5B",x"0C",x"17",x"2B",x"72",x"2B",x"73",x"D9",x"E5",x"D9",
x"D1",x"2B",x"72",x"2B",x"73",x"2B",x"36",x"2B",x"E5",x"FD",x"E1",x"C3",x"B1",x"DB",
x"FE",x"F5",x"D7",x"D9",x"2B",x"7E",x"FE",x"EC",x"20",x"FA",x"C3",x"A4",x"FF",x"08",
x"37",x"08",x"21",x"EB",x"E2",x"DD",x"36",x"05",x"20",x"37",x"D4",x"43",x"FC",x"FE",
x"BA",x"20",x"1F",x"CD",x"43",x"FC",x"CD",x"94",x"F2",x"FD",x"E5",x"CD",x"21",x"FA",
x"E1",x"23",x"D9",x"78",x"D9",x"08",x"B7",x"08",x"FE",x"A4",x"28",x"E2",x"FE",x"FD",
x"28",x"0C",x"30",x"0D",x"CF",x"01",x"CD",x"FB",x"FB",x"28",x"EC",x"08",x"30",x"F6",
x"D4",x"43",x"FC",x"3A",x"05",x"17",x"FE",x"20",x"CC",x"7F",x"FE",x"F7",x"24",x"CD",
x"4F",x"FF",x"20",x"A8",x"23",x"22",x"16",x"17",x"F6",x"37",x"08",x"D9",x"78",x"D9",
x"37",x"D4",x"43",x"FC",x"FE",x"FD",x"D2",x"B4",x"DB",x"E6",x"81",x"FE",x"01",x"C2",
x"5A",x"FD",x"08",x"30",x"49",x"2A",x"14",x"17",x"7D",x"B4",x"28",x"2E",x"7E",x"23",
x"FE",x"20",x"28",x"FA",x"2B",x"FE",x"21",x"28",x"19",x"FE",x"FD",x"38",x"33",x"D9",
x"E5",x"D5",x"C5",x"CD",x"C5",x"FC",x"D9",x"C1",x"D1",x"E1",x"D9",x"23",x"FE",x"FB",
x"28",x"E0",x"FE",x"FE",x"38",x"EB",x"2A",x"12",x"17",x"5E",x"16",x"00",x"19",x"22",
x"12",x"17",x"2A",x"12",x"17",x"7E",x"B7",x"28",x"0B",x"23",x"23",x"23",x"7E",x"23",
x"FE",x"20",x"28",x"FA",x"18",x"DC",x"CF",x"07",x"08",x"E5",x"D9",x"C5",x"CD",x"2F",
x"F4",x"C1",x"CB",x"49",x"E3",x"20",x"0B",x"CD",x"A1",x"F8",x"E3",x"CD",x"41",x"FB",
x"18",x"1E",x"CF",x"0C",x"CD",x"8E",x"FC",x"CD",x"14",x"F9",x"08",x"30",x"09",x"08",
x"30",x"F2",x"17",x"DA",x"12",x"F9",x"18",x"06",x"08",x"E5",x"CD",x"7F",x"EC",x"E1",
x"E3",x"CD",x"28",x"FB",x"E1",x"08",x"30",x"1A",x"08",x"7E",x"23",x"FE",x"20",x"28",
x"FA",x"FE",x"2C",x"28",x"0A",x"2B",x"FE",x"21",x"28",x"05",x"CB",x"7E",x"CA",x"92",
x"E2",x"22",x"14",x"17",x"18",x"0E",x"08",x"7E",x"23",x"FE",x"2C",x"28",x"04",x"3C",
x"20",x"F7",x"2B",x"22",x"16",x"17",x"D9",x"78",x"D9",x"FE",x"FD",x"D2",x"B4",x"DB",
x"FE",x"A4",x"CA",x"21",x"E2",x"CF",x"01",x"02",x"3F",x"20",x"DD",x"CB",x"02",x"C6",
x"CD",x"A7",x"F0",x"FD",x"7E",x"06",x"B7",x"08",x"CD",x"1B",x"FA",x"D9",x"E5",x"D9",
x"E1",x"3E",x"B5",x"CD",x"54",x"FD",x"08",x"28",x"13",x"08",x"18",x"08",x"23",x"E5",
x"D9",x"E1",x"D9",x"CD",x"43",x"FC",x"FE",x"02",x"CA",x"B2",x"E3",x"C3",x"81",x"DB",
x"FD",x"2A",x"1A",x"17",x"CD",x"C5",x"FC",x"FE",x"F4",x"28",x"E5",x"FE",x"FE",x"D2",
x"BB",x"DB",x"E5",x"D9",x"E1",x"D9",x"18",x"EE",x"DD",x"CB",x"02",x"C6",x"CD",x"1B",
x"FB",x"47",x"D9",x"78",x"D9",x"FE",x"EF",x"28",x"6E",x"FE",x"F0",x"20",x"24",x"CD",
x"57",x"E3",x"CD",x"DE",x"FB",x"FD",x"2A",x"1A",x"17",x"E5",x"CD",x"D1",x"FC",x"EB",
x"E1",x"18",x"37",x"CD",x"43",x"FC",x"05",x"C8",x"D9",x"E5",x"D9",x"E1",x"CD",x"43",
x"FC",x"30",x"06",x"FE",x"A4",x"28",x"EE",x"CF",x"01",x"D1",x"FD",x"2A",x"1A",x"17",
x"D9",x"CD",x"C5",x"FC",x"FE",x"F4",x"28",x"94",x"FE",x"FE",x"D2",x"14",x"FB",x"E5",
x"D9",x"E1",x"18",x"EE",x"CD",x"DE",x"FB",x"CD",x"43",x"FC",x"38",x"DF",x"D9",x"E5",
x"D9",x"D1",x"E5",x"CD",x"8E",x"FC",x"FD",x"E5",x"E1",x"2B",x"3A",x"02",x"17",x"77",
x"ED",x"4B",x"0C",x"17",x"2B",x"70",x"2B",x"71",x"2B",x"72",x"2B",x"73",x"2B",x"36",
x"06",x"E5",x"FD",x"E1",x"E1",x"18",x"0A",x"CD",x"57",x"E3",x"CD",x"DE",x"FB",x"FD",
x"2A",x"1A",x"17",x"C3",x"29",x"DE",x"2B",x"D9",x"CD",x"43",x"FC",x"E6",x"FD",x"FE",
x"01",x"C2",x"5A",x"FD",x"D9",x"CB",x"51",x"C2",x"5A",x"FD",x"CB",x"59",x"C4",x"0B",
x"F4",x"DD",x"71",x"01",x"D9",x"CD",x"2E",x"F4",x"D9",x"78",x"D9",x"E5",x"CD",x"E8",
x"E3",x"E1",x"CD",x"3B",x"FB",x"C3",x"B1",x"DB",x"D6",x"96",x"20",x"5E",x"CB",x"49",
x"C2",x"5A",x"FD",x"23",x"E5",x"4E",x"47",x"CD",x"27",x"FD",x"7A",x"BB",x"30",x"02",
x"7B",x"3D",x"57",x"79",x"92",x"E1",x"FD",x"E5",x"E5",x"D5",x"C5",x"38",x"0E",x"28",
x"0C",x"09",x"4F",x"FD",x"E5",x"D1",x"1B",x"ED",x"B8",x"13",x"D5",x"FD",x"E1",x"CD",
x"4A",x"E4",x"C1",x"D1",x"E1",x"7B",x"FD",x"E5",x"D1",x"13",x"FE",x"02",x"38",x"0C",
x"3D",x"B9",x"30",x"01",x"4F",x"09",x"0C",x"0D",x"28",x"02",x"ED",x"B8",x"E1",x"2B",
x"B7",x"ED",x"52",x"24",x"25",x"C2",x"12",x"F9",x"2C",x"CA",x"12",x"F9",x"2D",x"EB",
x"73",x"2B",x"36",x"01",x"E5",x"FD",x"E1",x"C9",x"3E",x"9A",x"CD",x"54",x"FD",x"C3",
x"8D",x"F2",x"CD",x"C4",x"FA",x"ED",x"5B",x"20",x"17",x"B7",x"ED",x"52",x"19",x"DA",
x"14",x"FB",x"ED",x"5B",x"22",x"17",x"ED",x"52",x"CA",x"B4",x"DB",x"E5",x"DC",x"86",
x"FC",x"4D",x"44",x"EB",x"38",x"13",x"D1",x"D5",x"E5",x"14",x"CA",x"14",x"FB",x"CD",
x"99",x"FC",x"E1",x"E5",x"CD",x"C9",x"DC",x"E1",x"09",x"18",x"08",x"B7",x"ED",x"42",
x"E5",x"CD",x"E9",x"DC",x"E1",x"22",x"22",x"17",x"C1",x"DD",x"CB",x"00",x"56",x"28",
x"0C",x"2A",x"0C",x"17",x"09",x"22",x"0C",x"17",x"C5",x"D9",x"D1",x"19",x"D9",x"CD",
x"FC",x"DC",x"C3",x"B1",x"DB",x"CF",x"08",x"D9",x"78",x"D9",x"FE",x"A4",x"C2",x"B4",
x"DB",x"CD",x"43",x"FC",x"DD",x"CB",x"00",x"D6",x"30",x"27",x"FE",x"03",x"28",x"07",
x"E6",x"82",x"C2",x"5A",x"FD",x"CF",x"0E",x"CD",x"2E",x"F4",x"EB",x"21",x"FD",x"09",
x"3E",x"2B",x"CD",x"E7",x"FC",x"38",x"D4",x"0E",x"05",x"09",x"0E",x"2B",x"7E",x"BB",
x"20",x"EE",x"23",x"7E",x"BA",x"20",x"E9",x"3E",x"2B",x"CD",x"E7",x"FC",x"38",x"BF",
x"23",x"5E",x"23",x"56",x"D5",x"23",x"5E",x"23",x"56",x"D5",x"23",x"5E",x"23",x"56",
x"D5",x"23",x"EB",x"11",x"22",x"00",x"FD",x"19",x"CD",x"63",x"FA",x"1B",x"21",x"F7",
x"FF",x"19",x"01",x"09",x"00",x"ED",x"B8",x"13",x"D5",x"FD",x"E1",x"FD",x"CB",x"08",
x"7E",x"F5",x"CD",x"93",x"F4",x"F1",x"E1",x"F5",x"FD",x"E5",x"CD",x"28",x"FB",x"FD",
x"E1",x"CD",x"93",x"F6",x"C1",x"D1",x"E1",x"79",x"17",x"30",x"06",x"28",x"07",x"F2",
x"AB",x"E4",x"AF",x"FA",x"AB",x"E4",x"ED",x"53",x"0C",x"17",x"11",x"D5",x"FF",x"FD",
x"19",x"C3",x"81",x"DB",x"CD",x"1B",x"FB",x"4F",x"3E",x"A4",x"CD",x"54",x"FD",x"CD",
x"1B",x"FB",x"ED",x"79",x"C3",x"B1",x"DB",x"CD",x"FF",x"FC",x"3E",x"A4",x"CD",x"54",
x"FD",x"CD",x"1B",x"FB",x"4F",x"CD",x"E7",x"FF",x"38",x"03",x"F3",x"D3",x"02",x"71",
x"3E",x"70",x"D3",x"02",x"FB",x"C3",x"B1",x"DB",x"0E",x"40",x"11",x"0E",x"20",x"DD",
x"71",x"05",x"08",x"AF",x"08",x"37",x"D4",x"43",x"FC",x"FE",x"AF",x"20",x"23",x"CD",
x"43",x"FC",x"CD",x"94",x"F2",x"21",x"31",x"18",x"36",x"7F",x"E5",x"CD",x"41",x"FB",
x"E1",x"23",x"5E",x"16",x"00",x"23",x"22",x"2E",x"17",x"19",x"72",x"22",x"30",x"17",
x"08",x"CB",x"C7",x"08",x"18",x"14",x"FE",x"B0",x"20",x"22",x"CD",x"16",x"FB",x"4F",
x"3E",x"A4",x"CD",x"54",x"FD",x"CD",x"1B",x"FB",x"47",x"CD",x"8B",x"E6",x"D9",x"78",
x"D9",x"08",x"B7",x"08",x"FE",x"A4",x"28",x"B8",x"FE",x"FD",x"28",x"0E",x"30",x"0F",
x"CF",x"01",x"CD",x"00",x"FC",x"28",x"EC",x"08",x"38",x"F6",x"08",x"37",x"D4",x"43",
x"FC",x"08",x"37",x"08",x"08",x"CB",x"47",x"F5",x"C4",x"9C",x"E6",x"F1",x"08",x"D9",
x"78",x"D9",x"FE",x"A4",x"20",x"06",x"3E",x"09",x"CD",x"9A",x"FE",x"C2",x"FE",x"A0",
x"20",x"08",x"CD",x"43",x"FC",x"08",x"B7",x"C3",x"7F",x"E6",x"FE",x"B6",x"20",x"15",
x"3E",x"96",x"CD",x"51",x"FD",x"CD",x"1B",x"FB",x"47",x"3E",x"95",x"CD",x"54",x"FD",
x"0E",x"00",x"CD",x"8B",x"E6",x"18",x"66",x"FE",x"FD",x"30",x"68",x"08",x"CB",x"47",
x"F5",x"28",x"17",x"08",x"2A",x"2E",x"17",x"ED",x"5B",x"30",x"17",x"B7",x"ED",x"52",
x"38",x"0B",x"21",x"33",x"18",x"22",x"2E",x"17",x"CD",x"9C",x"E6",x"08",x"08",x"D9",
x"78",x"D9",x"FE",x"02",x"30",x"25",x"CD",x"94",x"F2",x"17",x"30",x"23",x"F1",x"21",
x"9C",x"FF",x"C2",x"F0",x"FF",x"F6",x"FF",x"FD",x"E5",x"E1",x"23",x"F5",x"CD",x"7F",
x"FE",x"CD",x"21",x"FA",x"F1",x"3D",x"FA",x"7D",x"E6",x"F5",x"CD",x"C7",x"FE",x"18",
x"F5",x"CD",x"A7",x"F0",x"17",x"D2",x"5A",x"FD",x"F1",x"21",x"B5",x"FC",x"C2",x"F0",
x"FF",x"FD",x"E5",x"E1",x"23",x"CD",x"BA",x"FE",x"CD",x"1B",x"FA",x"08",x"37",x"08",
x"C3",x"DC",x"E5",x"08",x"DC",x"93",x"FE",x"08",x"C3",x"B4",x"DB",x"3A",x"05",x"17",
x"FE",x"20",x"28",x"03",x"FE",x"00",x"C0",x"F6",x"03",x"CD",x"1B",x"00",x"D7",x"C9",
x"ED",x"5B",x"30",x"17",x"2A",x"2E",x"17",x"7E",x"B7",x"ED",x"52",x"D0",x"19",x"E5",
x"21",x"BD",x"E6",x"01",x"0A",x"00",x"ED",x"B1",x"E1",x"C8",x"CD",x"9A",x"FE",x"23",
x"22",x"2E",x"17",x"18",x"E6",x"3C",x"3E",x"23",x"2A",x"25",x"2B",x"2D",x"24",x"5E",
x"2E",x"ED",x"5F",x"32",x"09",x"17",x"2A",x"1D",x"0B",x"22",x"0A",x"17",x"CD",x"D8",
x"E6",x"C3",x"B1",x"DB",x"06",x"10",x"3A",x"09",x"17",x"2A",x"0A",x"17",x"4F",x"0F",
x"0F",x"0F",x"A9",x"17",x"17",x"ED",x"6A",x"79",x"8F",x"10",x"F3",x"22",x"0A",x"17",
x"32",x"09",x"17",x"C9",x"2A",x"22",x"17",x"FE",x"02",x"20",x"06",x"CD",x"DE",x"FB",
x"CD",x"43",x"FC",x"22",x"12",x"17",x"21",x"00",x"00",x"22",x"14",x"17",x"C3",x"B4",
x"DB",x"CF",x"09",x"3E",x"06",x"CD",x"E7",x"FC",x"38",x"F7",x"DD",x"CB",x"00",x"D6",
x"23",x"5E",x"23",x"56",x"23",x"4E",x"23",x"46",x"ED",x"43",x"0C",x"17",x"23",x"7E",
x"32",x"02",x"17",x"23",x"E5",x"FD",x"E1",x"EB",x"C3",x"81",x"DB",x"CD",x"1B",x"FB",
x"0E",x"00",x"FE",x"02",x"28",x"0B",x"0C",x"FE",x"04",x"28",x"06",x"0C",x"FE",x"10",
x"C2",x"14",x"FB",x"F7",x"04",x"D7",x"C3",x"B1",x"DB",x"F7",x"08",x"CD",x"43",x"FC",
x"30",x"39",x"30",x"2C",x"FE",x"BE",x"20",x"05",x"F7",x"0A",x"D7",x"18",x"1B",x"FE",
x"A0",x"28",x"EA",x"FE",x"A4",x"28",x"1D",x"CD",x"C4",x"FA",x"4D",x"44",x"3E",x"A4",
x"CD",x"54",x"FD",x"CD",x"C4",x"FA",x"EB",x"F5",x"F7",x"06",x"D7",x"F1",x"FE",x"A0",
x"28",x"CF",x"FE",x"A4",x"28",x"02",x"F7",x"08",x"F7",x"09",x"D9",x"78",x"D9",x"FE",
x"FD",x"38",x"C2",x"C3",x"B4",x"DB",x"21",x"E4",x"E7",x"CD",x"12",x"FD",x"38",x"42",
x"CD",x"1B",x"FB",x"1E",x"00",x"32",x"1F",x"00",x"21",x"41",x"19",x"E5",x"06",x"7F",
x"1D",x"F2",x"B4",x"E7",x"D9",x"78",x"D9",x"FE",x"A4",x"20",x"1C",x"CD",x"43",x"FC",
x"FE",x"02",x"30",x"0D",x"CD",x"94",x"F2",x"21",x"3F",x"19",x"36",x"7F",x"CD",x"41",
x"FB",x"18",x"0D",x"CD",x"1B",x"FB",x"77",x"23",x"10",x"DA",x"04",x"36",x"00",x"23",
x"10",x"FB",x"D1",x"CD",x"1E",x"00",x"D7",x"D9",x"78",x"D9",x"FE",x"A0",x"C2",x"B4",
x"DB",x"CD",x"43",x"FC",x"18",x"AC",x"C3",x"11",x"B7",x"12",x"C4",x"13",x"BC",x"14",
x"C7",x"15",x"B9",x"16",x"C8",x"24",x"BD",x"2D",x"AE",x"34",x"00",x"1E",x"00",x"21",
x"1E",x"01",x"21",x"1E",x"02",x"21",x"1E",x"03",x"21",x"1E",x"1A",x"21",x"1E",x"1C",
x"16",x"00",x"21",x"4B",x"0B",x"19",x"CD",x"1B",x"FB",x"77",x"D9",x"78",x"D9",x"C9",
x"E1",x"E1",x"CD",x"1B",x"FB",x"4F",x"3E",x"0B",x"C3",x"9B",x"E7",x"E1",x"E1",x"3E",
x"0C",x"1E",x"01",x"C3",x"9D",x"E7",x"CD",x"1B",x"FB",x"87",x"32",x"4F",x"0B",x"18",
x"DF",x"21",x"15",x"0D",x"22",x"2A",x"17",x"21",x"07",x"32",x"22",x"2C",x"00",x"21",
x"15",x"0B",x"36",x"FF",x"37",x"D4",x"43",x"FC",x"FE",x"A0",x"28",x"23",x"21",x"7B",
x"E8",x"CD",x"12",x"FD",x"FE",x"A4",x"28",x"EF",x"F5",x"ED",x"5B",x"2A",x"17",x"ED",
x"4B",x"2C",x"00",x"F7",x"33",x"AF",x"32",x"15",x"0B",x"F1",x"FE",x"FD",x"30",x"0E",
x"FE",x"A0",x"C2",x"5A",x"FD",x"AF",x"32",x"15",x"0B",x"CD",x"43",x"FC",x"38",x"CD",
x"C3",x"B4",x"DB",x"BB",x"05",x"C6",x"0C",x"B3",x"0B",x"00",x"CD",x"C4",x"FA",x"22",
x"2A",x"17",x"F0",x"CF",x"04",x"F6",x"37",x"11",x"2C",x"00",x"38",x"01",x"13",x"CD",
x"1B",x"FB",x"12",x"D9",x"78",x"D9",x"C9",x"0E",x"50",x"CD",x"EE",x"FB",x"FE",x"E1",
x"28",x"0B",x"CB",x"F9",x"FE",x"FD",x"30",x"08",x"FE",x"EC",x"C2",x"5A",x"FD",x"CD",
x"43",x"FC",x"79",x"E6",x"7F",x"FE",x"50",x"28",x"04",x"FE",x"60",x"20",x"0A",x"79",
x"F6",x"04",x"CD",x"1B",x"00",x"D7",x"C3",x"B1",x"DB",x"CF",x"FF",x"0E",x"50",x"CD",
x"EE",x"FB",x"08",x"79",x"FE",x"50",x"28",x"04",x"FE",x"60",x"20",x"EF",x"F6",x"03",
x"4F",x"08",x"11",x"CE",x"19",x"FE",x"E1",x"28",x"0F",x"CB",x"F9",x"FE",x"02",x"38",
x"10",x"FE",x"FD",x"30",x"18",x"FE",x"EC",x"C2",x"5A",x"FD",x"CD",x"43",x"FC",x"FE",
x"02",x"30",x"0C",x"C5",x"CD",x"94",x"F2",x"FD",x"E5",x"CD",x"21",x"FA",x"D1",x"13",
x"C1",x"79",x"32",x"6B",x"0B",x"CD",x"1B",x"00",x"D7",x"C3",x"B1",x"DB",x"0E",x"10",
x"CD",x"EE",x"FB",x"08",x"79",x"F6",x"81",x"CD",x"1B",x"00",x"FD",x"E5",x"E1",x"FE",
x"EC",x"28",x"06",x"B7",x"D7",x"2B",x"71",x"3C",x"0E",x"AF",x"2B",x"77",x"2B",x"36",
x"01",x"08",x"FE",x"FD",x"D2",x"B4",x"DB",x"E5",x"FD",x"E1",x"FE",x"01",x"20",x"03",
x"D9",x"CB",x"51",x"C2",x"5A",x"FD",x"CB",x"59",x"C4",x"0B",x"F4",x"D9",x"CD",x"2E",
x"F4",x"CD",x"41",x"FB",x"C3",x"B1",x"DB",x"CD",x"35",x"EA",x"CD",x"10",x"DE",x"E5",
x"ED",x"5B",x"E1",x"19",x"D5",x"CD",x"99",x"FC",x"C1",x"D1",x"D5",x"3A",x"05",x"17",
x"F6",x"82",x"CD",x"1B",x"00",x"F5",x"C4",x"10",x"DE",x"F1",x"D7",x"CD",x"FC",x"DC",
x"CD",x"5A",x"EA",x"E1",x"3A",x"E3",x"19",x"B7",x"CA",x"DA",x"DA",x"C3",x"23",x"DE",
x"AF",x"CD",x"FB",x"E9",x"11",x"EF",x"19",x"06",x"10",x"AF",x"1B",x"12",x"10",x"FC",
x"D5",x"3C",x"32",x"E0",x"19",x"3A",x"07",x"17",x"32",x"E3",x"19",x"CD",x"41",x"DD",
x"23",x"ED",x"5B",x"22",x"17",x"AF",x"32",x"07",x"17",x"ED",x"52",x"22",x"E1",x"19",
x"E3",x"D5",x"06",x"10",x"3A",x"05",x"17",x"F6",x"01",x"32",x"1F",x"00",x"4E",x"23",
x"C5",x"CD",x"1E",x"00",x"D7",x"C1",x"10",x"F6",x"D1",x"C1",x"3A",x"05",x"17",x"F6",
x"02",x"CD",x"1B",x"00",x"D7",x"CD",x"5A",x"EA",x"C3",x"B1",x"DB",x"CD",x"35",x"EA",
x"CD",x"41",x"DD",x"23",x"ED",x"5B",x"22",x"17",x"B7",x"ED",x"52",x"ED",x"4B",x"E1",
x"19",x"ED",x"42",x"C2",x"58",x"EA",x"3A",x"05",x"17",x"F6",x"85",x"CD",x"1B",x"00",
x"D7",x"CD",x"5A",x"EA",x"C3",x"B1",x"DB",x"3E",x"80",x"DD",x"CB",x"00",x"DE",x"F5",
x"0E",x"50",x"CD",x"EE",x"FB",x"08",x"79",x"FE",x"50",x"28",x"05",x"FE",x"60",x"C2",
x"C7",x"E8",x"C1",x"B0",x"32",x"05",x"17",x"F6",x"03",x"32",x"1F",x"00",x"08",x"11",
x"CE",x"19",x"FE",x"02",x"30",x"0A",x"CD",x"94",x"F2",x"FD",x"E5",x"CD",x"21",x"FA",
x"D1",x"13",x"AF",x"32",x"6B",x"0B",x"CD",x"1E",x"00",x"D7",x"C9",x"CD",x"F9",x"E9",
x"3A",x"05",x"17",x"F6",x"81",x"32",x"1F",x"00",x"21",x"DF",x"19",x"E5",x"06",x"10",
x"C5",x"CD",x"1E",x"00",x"D7",x"71",x"23",x"C1",x"10",x"F6",x"E1",x"B6",x"20",x"04",
x"23",x"3C",x"96",x"C8",x"CF",x"10",x"3A",x"05",x"17",x"F6",x"04",x"CD",x"1B",x"00",
x"D7",x"DD",x"CB",x"00",x"9E",x"C9",x"3E",x"96",x"CD",x"54",x"FD",x"CD",x"A7",x"F0",
x"3E",x"95",x"C3",x"54",x"FD",x"3E",x"96",x"CD",x"54",x"FD",x"CD",x"94",x"F2",x"3E",
x"95",x"C3",x"54",x"FD",x"2A",x"18",x"17",x"7E",x"23",x"22",x"18",x"17",x"6F",x"AF",
x"67",x"E5",x"29",x"29",x"29",x"D1",x"ED",x"52",x"11",x"11",x"C1",x"19",x"18",x"08",
x"21",x"C7",x"19",x"18",x"03",x"21",x"C0",x"19",x"CD",x"8E",x"FC",x"11",x"06",x"00",
x"19",x"FD",x"E5",x"D1",x"1B",x"ED",x"A8",x"AF",x"12",x"1B",x"01",x"06",x"00",x"ED",
x"B8",x"3E",x"09",x"12",x"D5",x"FD",x"E1",x"C9",x"11",x"C7",x"19",x"18",x"03",x"11",
x"C0",x"19",x"CD",x"D5",x"EA",x"E5",x"FD",x"E1",x"C9",x"11",x"C7",x"19",x"18",x"03",
x"11",x"C0",x"19",x"FD",x"E5",x"E1",x"23",x"01",x"06",x"00",x"ED",x"B0",x"23",x"ED",
x"A0",x"C9",x"00",x"00",x"03",x"41",x"42",x"53",x"0A",x"CD",x"68",x"EA",x"FD",x"CB",
x"08",x"BE",x"C9",x"CD",x"43",x"FC",x"CD",x"68",x"EA",x"01",x"00",x"00",x"FD",x"7E",
x"08",x"E6",x"80",x"4F",x"C5",x"C4",x"26",x"F7",x"DF",x"08",x"85",x"01",x"CD",x"93",
x"F6",x"FA",x"1A",x"EB",x"28",x"0A",x"C1",x"06",x"02",x"C5",x"DF",x"05",x"01",x"06",
x"01",x"8A",x"DF",x"06",x"85",x"02",x"CD",x"93",x"F6",x"FA",x"3C",x"EB",x"28",x"16",
x"C1",x"04",x"C5",x"DF",x"05",x"04",x"06",x"02",x"05",x"00",x"03",x"05",x"00",x"03",
x"06",x"00",x"05",x"03",x"06",x"00",x"01",x"8A",x"DF",x"06",x"0C",x"0C",x"0C",x"02",
x"08",x"05",x"06",x"02",x"05",x"05",x"00",x"06",x"02",x"06",x"05",x"08",x"00",x"06",
x"02",x"05",x"07",x"00",x"01",x"02",x"80",x"C1",x"78",x"FE",x"02",x"D4",x"26",x"F7",
x"C5",x"21",x"14",x"C2",x"05",x"28",x"0C",x"21",x"06",x"C2",x"05",x"28",x"06",x"21",
x"0D",x"C2",x"05",x"20",x"06",x"CD",x"A2",x"EA",x"CD",x"93",x"F4",x"C1",x"79",x"FD",
x"AE",x"08",x"FD",x"77",x"08",x"C9",x"E2",x"EA",x"04",x"43",x"48",x"52",x"24",x"08",
x"CD",x"68",x"EA",x"CD",x"1A",x"FB",x"FD",x"E5",x"E1",x"2B",x"77",x"2B",x"36",x"01",
x"2B",x"36",x"01",x"E5",x"FD",x"E1",x"C9",x"80",x"EB",x"03",x"43",x"4F",x"53",x"0A",
x"CD",x"68",x"EA",x"DF",x"05",x"23",x"80",x"C3",x"5E",x"EE",x"9D",x"EB",x"03",x"45",
x"58",x"50",x"0A",x"CD",x"68",x"EA",x"DF",x"0C",x"05",x"09",x"82",x"CD",x"AF",x"EC",
x"FD",x"7E",x"08",x"4F",x"E6",x"7F",x"FE",x"43",x"38",x"0A",x"B1",x"F2",x"12",x"F9",
x"CD",x"1B",x"FA",x"C3",x"F9",x"F9",x"CD",x"92",x"FA",x"CD",x"C3",x"FA",x"5D",x"54",
x"01",x"7E",x"00",x"B7",x"ED",x"4A",x"FA",x"CE",x"EB",x"CB",x"21",x"ED",x"42",x"D2",
x"12",x"F9",x"D5",x"DF",x"09",x"05",x"0A",x"02",x"03",x"07",x"05",x"0B",x"02",x"03",
x"0C",x"0C",x"02",x"08",x"05",x"10",x"00",x"06",x"02",x"05",x"0F",x"00",x"0B",x"05",
x"0E",x"06",x"02",x"05",x"0D",x"00",x"06",x"02",x"05",x"0C",x"00",x"02",x"08",x"07",
x"06",x"03",x"01",x"05",x"00",x"00",x"0C",x"00",x"8A",x"D1",x"CB",x"43",x"28",x"15",
x"D5",x"DF",x"06",x"05",x"20",x"02",x"8A",x"D1",x"14",x"15",x"13",x"28",x"08",x"FA",
x"37",x"EC",x"21",x"C6",x"19",x"34",x"1B",x"21",x"C6",x"19",x"AF",x"B3",x"1F",x"86",
x"E6",x"7F",x"77",x"C3",x"9F",x"EA",x"AE",x"EB",x"04",x"46",x"52",x"45",x"45",x"0A",
x"FD",x"E5",x"E1",x"ED",x"5B",x"26",x"17",x"B7",x"ED",x"52",x"11",x"00",x"01",x"ED",
x"52",x"11",x"FF",x"7F",x"ED",x"52",x"D5",x"CD",x"2B",x"FA",x"E1",x"CD",x"2B",x"FA",
x"C3",x"93",x"F4",x"44",x"EC",x"02",x"49",x"4E",x"0A",x"CD",x"68",x"EA",x"CD",x"1A",
x"FB",x"4F",x"ED",x"68",x"26",x"00",x"C3",x"2B",x"FA",x"D0",x"17",x"D0",x"CD",x"1B",
x"FA",x"DF",x"85",x"27",x"C9",x"CD",x"43",x"FC",x"F7",x"93",x"D7",x"FD",x"E5",x"E1",
x"2B",x"79",x"B7",x"28",x"06",x"F7",x"91",x"D7",x"71",x"2B",x"3C",x"77",x"2B",x"36",
x"01",x"E5",x"FD",x"E1",x"C9",x"6B",x"EC",x"03",x"49",x"4E",x"54",x"0A",x"CD",x"68",
x"EA",x"FD",x"7E",x"08",x"E6",x"7F",x"D6",x"40",x"38",x"20",x"3C",x"F5",x"CD",x"07",
x"F7",x"CD",x"DF",x"F9",x"F1",x"C6",x"03",x"47",x"3E",x"00",x"DC",x"E3",x"F7",x"04",
x"78",x"FE",x"10",x"38",x"F5",x"CD",x"07",x"F7",x"CD",x"DF",x"F9",x"C3",x"34",x"F7",
x"FD",x"7E",x"08",x"B7",x"F2",x"F9",x"F9",x"CD",x"08",x"FA",x"C3",x"26",x"F7",x"A5",
x"EC",x"02",x"49",x"4F",x"0A",x"CD",x"68",x"EA",x"CD",x"1A",x"FB",x"6F",x"26",x"00",
x"11",x"41",x"19",x"29",x"19",x"5E",x"23",x"56",x"EB",x"C3",x"2B",x"FA",x"E5",x"EC",
x"03",x"4C",x"45",x"4E",x"0A",x"CD",x"75",x"EA",x"FD",x"E5",x"CD",x"21",x"FA",x"E1",
x"23",x"6E",x"26",x"00",x"C3",x"2B",x"FA",x"00",x"ED",x"03",x"4C",x"4F",x"47",x"0A",
x"CD",x"68",x"EA",x"CD",x"C3",x"EA",x"21",x"C5",x"19",x"AF",x"57",x"B6",x"CA",x"14",
x"FB",x"23",x"5E",x"1C",x"1D",x"FA",x"14",x"FB",x"36",x"3F",x"D5",x"E5",x"DF",x"06",
x"85",x"20",x"CD",x"93",x"F6",x"E1",x"28",x"03",x"F2",x"49",x"ED",x"D1",x"1B",x"34",
x"D5",x"DF",x"06",x"05",x"00",x"03",x"05",x"00",x"03",x"06",x"05",x"01",x"00",x"01",
x"08",x"0C",x"0C",x"02",x"08",x"05",x"14",x"02",x"05",x"13",x"00",x"06",x"02",x"05",
x"12",x"00",x"06",x"02",x"06",x"05",x"17",x"00",x"06",x"02",x"05",x"16",x"00",x"06",
x"02",x"05",x"15",x"00",x"01",x"05",x"18",x"00",x"82",x"E1",x"11",x"3F",x"00",x"B7",
x"ED",x"52",x"CD",x"2B",x"FA",x"DF",x"00",x"05",x"11",x"82",x"C9",x"CD",x"A6",x"FA",
x"CD",x"D2",x"EA",x"CD",x"FB",x"F5",x"CD",x"AF",x"EC",x"DF",x"02",x"03",x"8C",x"FD",
x"CB",x"08",x"BE",x"CD",x"9F",x"EA",x"CD",x"93",x"F6",x"F8",x"C3",x"F9",x"F9",x"CD",
x"43",x"FC",x"CD",x"75",x"EA",x"FD",x"E5",x"CD",x"21",x"FA",x"E1",x"23",x"7E",x"B7",
x"CA",x"14",x"FB",x"C3",x"10",x"ED",x"17",x"ED",x"04",x"50",x"45",x"45",x"4B",x"0A",
x"CD",x"68",x"EA",x"CD",x"02",x"FD",x"CD",x"E7",x"FF",x"38",x"03",x"F3",x"D3",x"02",
x"6E",x"3E",x"70",x"D3",x"02",x"FB",x"C3",x"12",x"ED",x"BE",x"ED",x"02",x"50",x"49",
x"0A",x"DF",x"85",x"22",x"C9",x"DD",x"ED",x"03",x"52",x"4E",x"44",x"0A",x"FE",x"96",
x"28",x"10",x"CD",x"D8",x"E6",x"CD",x"2B",x"FA",x"DF",x"05",x"26",x"00",x"05",x"26",
x"0C",x"00",x"81",x"C9",x"CD",x"68",x"EA",x"CD",x"C3",x"FA",x"CB",x"7C",x"C2",x"14",
x"FB",x"7C",x"B5",x"CA",x"14",x"FB",x"E5",x"AF",x"3C",x"29",x"30",x"FC",x"3D",x"E1",
x"2B",x"E5",x"F5",x"CD",x"D8",x"E6",x"F1",x"47",x"CB",x"3C",x"CB",x"1D",x"10",x"FA",
x"EB",x"E1",x"B7",x"ED",x"52",x"19",x"38",x"EB",x"EB",x"C3",x"2B",x"FA",x"E7",x"ED",
x"03",x"53",x"47",x"4E",x"0A",x"CD",x"68",x"EA",x"FD",x"7E",x"06",x"B7",x"C8",x"FD",
x"7E",x"08",x"F5",x"CD",x"08",x"FA",x"F1",x"E6",x"80",x"FD",x"B6",x"08",x"FD",x"77",
x"08",x"C9",x"34",x"EE",x"03",x"53",x"49",x"4E",x"0A",x"CD",x"68",x"EA",x"DF",x"05",
x"22",x"05",x"22",x"80",x"CD",x"8B",x"ED",x"FD",x"7E",x"08",x"B7",x"1F",x"F5",x"DF",
x"8A",x"DF",x"06",x"85",x"23",x"F1",x"F5",x"FC",x"26",x"F7",x"CD",x"93",x"F6",x"C1",
x"C5",x"28",x"1B",x"A8",x"FA",x"93",x"EE",x"DF",x"06",x"85",x"22",x"F1",x"EE",x"40",
x"F5",x"F4",x"26",x"F7",x"DF",x"00",x"8A",x"18",x"DC",x"F1",x"EE",x"80",x"F5",x"FA",
x"6F",x"EE",x"DF",x"06",x"0C",x"0C",x"0C",x"02",x"08",x"05",x"1D",x"02",x"05",x"1C",
x"00",x"06",x"02",x"05",x"1B",x"00",x"06",x"02",x"05",x"1A",x"00",x"06",x"02",x"05",
x"19",x"00",x"06",x"02",x"02",x"80",x"F1",x"87",x"F0",x"C3",x"26",x"F7",x"54",x"EE",
x"03",x"53",x"51",x"52",x"0A",x"CD",x"68",x"EA",x"FD",x"CB",x"08",x"7E",x"C2",x"14",
x"FB",x"FD",x"7E",x"06",x"B7",x"C8",x"CD",x"C3",x"EA",x"21",x"C6",x"19",x"7E",x"D6",
x"3F",x"F5",x"36",x"3F",x"DF",x"06",x"05",x"1F",x"02",x"05",x"1E",x"00",x"8B",x"06",
x"04",x"C5",x"DF",x"07",x"06",x"07",x"01",x"07",x"03",x"05",x"00",x"02",x"00",x"8B",
x"C1",x"10",x"F0",x"F1",x"CB",x"47",x"28",x"09",x"F5",x"DF",x"07",x"05",x"20",x"02",
x"8B",x"F1",x"3C",x"CB",x"3F",x"21",x"CD",x"19",x"86",x"E6",x"7F",x"77",x"C3",x"9A",
x"EA",x"FD",x"7E",x"06",x"B7",x"20",x"06",x"CD",x"1B",x"FA",x"C3",x"08",x"FA",x"FD",
x"7E",x"0F",x"B7",x"CA",x"1B",x"FA",x"FD",x"7E",x"08",x"E6",x"7F",x"FE",x"43",x"30",
x"4A",x"CD",x"92",x"FA",x"CD",x"C3",x"FA",x"E5",x"CD",x"92",x"FA",x"CD",x"67",x"F7",
x"E1",x"E5",x"CD",x"2B",x"FA",x"CD",x"93",x"F6",x"E1",x"20",x"32",x"CB",x"7C",x"F5",
x"C4",x"86",x"FC",x"E5",x"DF",x"0A",x"0A",x"85",x"01",x"E1",x"E5",x"CB",x"45",x"28",
x"06",x"CD",x"9F",x"EA",x"CD",x"12",x"F5",x"E1",x"CB",x"3C",x"CB",x"1D",x"7C",x"B5",
x"28",x"08",x"E5",x"DF",x"06",x"06",x"02",x"8A",x"18",x"E3",x"F1",x"C8",x"DF",x"0B",
x"05",x"01",x"07",x"81",x"C9",x"CD",x"BE",x"EA",x"CD",x"21",x"ED",x"CD",x"9A",x"EA",
x"CD",x"12",x"F5",x"C3",x"B8",x"EB",x"C0",x"EE",x"04",x"53",x"54",x"52",x"24",x"08",
x"CD",x"68",x"EA",x"CD",x"0E",x"F8",x"CD",x"1B",x"FA",x"C3",x"7D",x"FA",x"8C",x"EF",
x"07",x"53",x"54",x"52",x"49",x"4E",x"47",x"24",x"08",x"3E",x"96",x"CD",x"54",x"FD",
x"CD",x"1B",x"FB",x"F5",x"3E",x"A4",x"CD",x"54",x"FD",x"FE",x"02",x"30",x"13",x"CD",
x"94",x"F2",x"FD",x"7E",x"01",x"B7",x"28",x"07",x"FD",x"7E",x"02",x"CD",x"21",x"FA",
x"01",x"C1",x"F5",x"37",x"D4",x"1B",x"FB",x"F5",x"CD",x"70",x"EA",x"D1",x"FD",x"E5",
x"E1",x"2B",x"F1",x"3C",x"CA",x"12",x"F9",x"3D",x"28",x"05",x"47",x"72",x"2B",x"10",
x"FC",x"77",x"2B",x"36",x"01",x"E5",x"FD",x"E1",x"C9",x"A0",x"EF",x"03",x"54",x"41",
x"4E",x"0A",x"CD",x"68",x"EA",x"CD",x"CD",x"EA",x"CD",x"5E",x"EE",x"DF",x"07",x"05",
x"23",x"80",x"CD",x"5E",x"EE",x"C3",x"FB",x"F5",x"F1",x"EF",x"03",x"55",x"53",x"52",
x"0A",x"3E",x"96",x"CD",x"54",x"FD",x"CD",x"A7",x"F0",x"FE",x"95",x"28",x"0A",x"3E",
x"A4",x"CD",x"54",x"FD",x"CD",x"C4",x"FA",x"3E",x"95",x"CD",x"54",x"FD",x"11",x"2B",
x"FA",x"D5",x"E5",x"CD",x"02",x"FD",x"E3",x"C9",x"0C",x"F0",x"03",x"56",x"41",x"4C",
x"0A",x"CD",x"75",x"EA",x"FD",x"E5",x"E1",x"23",x"E5",x"4E",x"06",x"00",x"09",x"23",
x"7E",x"70",x"E3",x"F5",x"23",x"CD",x"14",x"F9",x"CD",x"7F",x"EC",x"F1",x"E1",x"77",
x"2B",x"EB",x"FD",x"E5",x"E1",x"01",x"09",x"00",x"09",x"2B",x"ED",x"B8",x"13",x"D5",
x"FD",x"E1",x"C9",x"36",x"F0",x"06",x"56",x"41",x"52",x"50",x"54",x"52",x"0A",x"3E",
x"96",x"CD",x"54",x"FD",x"E6",x"FD",x"FE",x"01",x"C2",x"14",x"FB",x"D9",x"79",x"E6",
x"7F",x"32",x"08",x"17",x"E6",x"0C",x"20",x"F2",x"D9",x"CD",x"2E",x"F4",x"CD",x"2B",
x"FA",x"C3",x"70",x"EA",x"69",x"F0",x"06",x"56",x"45",x"52",x"4E",x"55",x"4D",x"0A",
x"21",x"0C",x"00",x"C3",x"2B",x"FA",x"CD",x"43",x"FC",x"D9",x"78",x"D9",x"CD",x"D7",
x"F0",x"D9",x"78",x"D9",x"FE",x"BF",x"28",x"04",x"FE",x"B2",x"C0",x"37",x"F5",x"CD",
x"43",x"FC",x"CD",x"D7",x"F0",x"CD",x"BF",x"FA",x"F1",x"38",x"07",x"7D",x"B3",x"6F",
x"7C",x"B2",x"18",x"05",x"7D",x"AB",x"6F",x"7C",x"B2",x"67",x"CD",x"2B",x"FA",x"18",
x"D6",x"CD",x"F4",x"F0",x"D9",x"78",x"D9",x"FE",x"C9",x"C0",x"CD",x"43",x"FC",x"CD",
x"F4",x"F0",x"CD",x"BF",x"FA",x"7D",x"A3",x"6F",x"7C",x"A2",x"67",x"CD",x"2B",x"FA",
x"18",x"E6",x"FE",x"C2",x"20",x"12",x"CD",x"43",x"FC",x"CD",x"F4",x"F0",x"CD",x"C3",
x"FA",x"7D",x"2F",x"6F",x"7C",x"2F",x"67",x"C3",x"2B",x"FA",x"FE",x"02",x"38",x"15",
x"CD",x"55",x"F1",x"FE",x"99",x"D8",x"FE",x"9F",x"D0",x"F5",x"CD",x"43",x"FC",x"CD",
x"55",x"F1",x"CD",x"93",x"F6",x"18",x"17",x"CD",x"94",x"F2",x"FE",x"99",x"DA",x"5D",
x"F3",x"FE",x"9F",x"D2",x"5D",x"F3",x"F5",x"CD",x"43",x"FC",x"CD",x"94",x"F2",x"CD",
x"D7",x"F6",x"E1",x"7C",x"CD",x"42",x"F1",x"C3",x"2B",x"FA",x"21",x"FF",x"FF",x"0F",
x"30",x"01",x"F8",x"0F",x"30",x"01",x"C8",x"0F",x"30",x"03",x"28",x"01",x"F0",x"23",
x"C9",x"CD",x"6C",x"F1",x"C4",x"81",x"F1",x"1C",x"C4",x"26",x"F7",x"CD",x"6C",x"F1",
x"C0",x"1C",x"CC",x"93",x"F4",x"C4",x"8E",x"F4",x"18",x"F3",x"D9",x"78",x"D9",x"1E",
x"FF",x"FE",x"98",x"28",x"04",x"FE",x"A2",x"C0",x"1C",x"CD",x"43",x"FC",x"CD",x"81",
x"F1",x"AF",x"C9",x"CD",x"A2",x"F1",x"D9",x"78",x"D9",x"FE",x"A8",x"28",x"03",x"FE",
x"A1",x"C0",x"57",x"CD",x"43",x"FC",x"CD",x"A2",x"F1",x"D5",x"7A",x"FE",x"A8",x"CC",
x"12",x"F5",x"C4",x"FB",x"F5",x"D1",x"18",x"E2",x"D5",x"CD",x"BB",x"F1",x"D1",x"D9",
x"78",x"D9",x"FE",x"9F",x"C0",x"D5",x"CD",x"43",x"FC",x"CD",x"BB",x"F1",x"CD",x"17",
x"EF",x"18",x"ED",x"CF",x"03",x"F5",x"CD",x"8E",x"FC",x"F1",x"FE",x"C0",x"CA",x"A9",
x"ED",x"FE",x"B1",x"CA",x"F1",x"EA",x"FE",x"02",x"DA",x"5D",x"F3",x"CA",x"43",x"FC",
x"FE",x"FD",x"30",x"E3",x"FE",x"96",x"20",x"08",x"CD",x"A4",x"F0",x"FE",x"95",x"CA",
x"43",x"FC",x"FE",x"03",x"C2",x"5A",x"FD",x"CD",x"2E",x"F4",x"CB",x"59",x"C2",x"AD",
x"DB",x"CB",x"51",x"CA",x"63",x"FA",x"DD",x"56",x"01",x"D5",x"E5",x"D6",x"96",x"D6",
x"01",x"9F",x"F5",x"79",x"28",x"14",x"08",x"CD",x"43",x"FC",x"B7",x"FA",x"5A",x"FD",
x"DD",x"77",x"01",x"CD",x"8D",x"F2",x"3E",x"95",x"CD",x"54",x"FD",x"08",x"08",x"F1",
x"2A",x"26",x"17",x"E3",x"E5",x"2A",x"24",x"17",x"E3",x"D9",x"E5",x"2A",x"0C",x"17",
x"E5",x"C5",x"D9",x"5E",x"23",x"56",x"23",x"ED",x"53",x"0C",x"17",x"5E",x"23",x"56",
x"EB",x"D9",x"4F",x"CD",x"43",x"FC",x"D6",x"96",x"D6",x"01",x"9F",x"A9",x"C2",x"5A",
x"FD",x"A9",x"28",x"27",x"CD",x"43",x"FC",x"E6",x"81",x"FE",x"01",x"C2",x"5A",x"FD",
x"D9",x"CB",x"79",x"CC",x"0B",x"F4",x"79",x"DD",x"AE",x"01",x"E6",x"02",x"C2",x"5D",
x"F3",x"D5",x"D9",x"E1",x"CD",x"3B",x"FB",x"CD",x"43",x"FC",x"3E",x"95",x"CD",x"54",
x"FD",x"3E",x"9A",x"CD",x"54",x"FD",x"08",x"DD",x"77",x"01",x"CD",x"8D",x"F2",x"C1",
x"E1",x"22",x"0C",x"17",x"E1",x"D9",x"E1",x"22",x"24",x"17",x"E1",x"22",x"26",x"17",
x"F1",x"32",x"01",x"17",x"C9",x"DD",x"CB",x"01",x"4E",x"C2",x"A7",x"F0",x"D9",x"78",
x"D9",x"CD",x"E0",x"F2",x"D9",x"78",x"D9",x"FE",x"97",x"C0",x"CD",x"43",x"FC",x"CD",
x"E0",x"F2",x"FD",x"E5",x"E1",x"23",x"5D",x"54",x"4E",x"06",x"00",x"09",x"23",x"E5",
x"FD",x"E1",x"23",x"4E",x"CD",x"8E",x"FC",x"E5",x"09",x"79",x"B7",x"1A",x"28",x"02",
x"ED",x"B8",x"E1",x"86",x"12",x"DA",x"12",x"F9",x"FE",x"FF",x"CA",x"12",x"F9",x"4E",
x"5D",x"54",x"1B",x"1B",x"09",x"EB",x"4F",x"03",x"ED",x"B8",x"EB",x"36",x"01",x"E5",
x"FD",x"E1",x"18",x"BA",x"CD",x"2D",x"F3",x"D9",x"78",x"D9",x"FE",x"96",x"C0",x"CD",
x"27",x"FD",x"FD",x"E5",x"E1",x"23",x"7E",x"4F",x"06",x"00",x"BA",x"38",x"01",x"7A",
x"57",x"B7",x"28",x"0D",x"79",x"BB",x"38",x"09",x"1C",x"1D",x"20",x"01",x"1C",x"7A",
x"93",x"30",x"04",x"09",x"AF",x"18",x"0B",x"3C",x"E5",x"09",x"EB",x"4C",x"E1",x"09",
x"4F",x"ED",x"B8",x"EB",x"77",x"2B",x"36",x"01",x"E5",x"FD",x"E1",x"18",x"C2",x"CD",
x"C4",x"FA",x"16",x"00",x"24",x"C8",x"15",x"25",x"C0",x"55",x"C9",x"CD",x"8E",x"FC",
x"D9",x"C5",x"D9",x"C1",x"78",x"FE",x"01",x"DA",x"43",x"FC",x"28",x"0B",x"FE",x"04",
x"38",x"1D",x"FE",x"FD",x"DA",x"5A",x"FD",x"CF",x"03",x"79",x"FE",x"C5",x"CA",x"89",
x"EC",x"CD",x"2E",x"F4",x"CB",x"59",x"C2",x"AD",x"DB",x"CB",x"51",x"C2",x"F4",x"F1",
x"C3",x"7C",x"FA",x"CF",x"0E",x"CD",x"8E",x"FC",x"ED",x"5B",x"24",x"17",x"2A",x"26",
x"17",x"22",x"24",x"17",x"73",x"23",x"72",x"23",x"0E",x"00",x"E5",x"ED",x"5B",x"28",
x"17",x"1A",x"FE",x"FD",x"30",x"27",x"FE",x"20",x"38",x"1C",x"FE",x"24",x"28",x"19",
x"FE",x"2E",x"28",x"14",x"FE",x"30",x"38",x"17",x"FE",x"3A",x"38",x"0C",x"FE",x"3F",
x"38",x"0F",x"FE",x"60",x"38",x"04",x"FE",x"A9",x"38",x"07",x"37",x"13",x"0C",x"23",
x"77",x"38",x"D4",x"7E",x"23",x"22",x"26",x"17",x"E3",x"71",x"E1",x"C9",x"CD",x"8E",
x"FC",x"2A",x"26",x"17",x"06",x"06",x"AF",x"77",x"23",x"10",x"FC",x"18",x"13",x"DD",
x"CB",x"01",x"4E",x"20",x"EB",x"CD",x"8E",x"FC",x"2A",x"26",x"17",x"71",x"23",x"06",
x"00",x"70",x"09",x"23",x"22",x"26",x"17",x"C9",x"22",x"28",x"17",x"21",x"25",x"17",
x"3E",x"E1",x"56",x"2B",x"5E",x"7B",x"B2",x"2A",x"28",x"17",x"C8",x"EB",x"23",x"E5",
x"23",x"46",x"1A",x"13",x"23",x"BE",x"20",x"EB",x"10",x"F8",x"FE",x"24",x"28",x"10",
x"1A",x"FE",x"20",x"28",x"0B",x"FE",x"FD",x"30",x"07",x"FE",x"A9",x"30",x"D8",x"17",
x"30",x"D5",x"F1",x"23",x"CB",x"BE",x"37",x"18",x"1D",x"CD",x"5F",x"F3",x"D6",x"24",
x"28",x"02",x"3E",x"02",x"77",x"E5",x"23",x"22",x"26",x"17",x"20",x"06",x"0E",x"12",
x"CD",x"C1",x"F3",x"AF",x"C4",x"AC",x"F3",x"E1",x"CB",x"FE",x"4E",x"23",x"EB",x"C9",
x"CF",x"05",x"D9",x"D5",x"CB",x"41",x"79",x"D9",x"E1",x"4F",x"CA",x"43",x"FC",x"3E",
x"96",x"CD",x"51",x"FD",x"AF",x"5F",x"57",x"7E",x"23",x"EB",x"C5",x"E5",x"F5",x"3E",
x"A4",x"C4",x"54",x"FD",x"CD",x"C4",x"FA",x"EB",x"4E",x"23",x"46",x"23",x"EB",x"B7",
x"ED",x"42",x"30",x"D2",x"09",x"F1",x"F5",x"D5",x"3D",x"28",x"0E",x"EB",x"4E",x"23",
x"46",x"23",x"E5",x"F5",x"CD",x"B3",x"FC",x"F1",x"D1",x"18",x"EF",x"D1",x"F1",x"C1",
x"09",x"3D",x"20",x"CF",x"3E",x"95",x"CD",x"54",x"FD",x"EB",x"C1",x"CB",x"49",x"01",
x"06",x"00",x"20",x"03",x"4E",x"03",x"03",x"E5",x"CD",x"B3",x"FC",x"D1",x"19",x"C9",
x"F5",x"CD",x"26",x"F7",x"F1",x"F5",x"FD",x"E5",x"11",x"09",x"00",x"FD",x"19",x"FD",
x"E3",x"FD",x"7E",x"08",x"E6",x"7F",x"4F",x"FD",x"7E",x"11",x"E6",x"7F",x"91",x"F2",
x"BF",x"F4",x"FD",x"E3",x"F5",x"ED",x"44",x"CD",x"90",x"F7",x"C1",x"FD",x"E3",x"FD",
x"7E",x"11",x"90",x"FD",x"77",x"11",x"AF",x"C4",x"90",x"F7",x"FD",x"7E",x"08",x"FD",
x"AE",x"11",x"07",x"D4",x"F4",x"F4",x"FD",x"E3",x"30",x"1E",x"CD",x"1C",x"F7",x"FD",
x"E3",x"CD",x"1C",x"F7",x"CD",x"F4",x"F4",x"FD",x"E3",x"FD",x"7E",x"07",x"B7",x"28",
x"0B",x"CD",x"0C",x"F7",x"3E",x"80",x"FD",x"AE",x"08",x"FD",x"77",x"08",x"F1",x"CD",
x"34",x"F7",x"F1",x"C9",x"F5",x"FD",x"E5",x"D1",x"21",x"09",x"00",x"19",x"06",x"07",
x"23",x"13",x"1A",x"8E",x"27",x"77",x"10",x"F8",x"F1",x"C9",x"11",x"09",x"00",x"FD",
x"19",x"CD",x"F9",x"F9",x"F1",x"C9",x"F5",x"FD",x"7E",x"0F",x"B7",x"28",x"EF",x"FD",
x"7E",x"06",x"B7",x"28",x"E9",x"FD",x"7E",x"11",x"FD",x"6E",x"08",x"AD",x"67",x"AD",
x"E6",x"7F",x"6F",x"FD",x"7E",x"08",x"E6",x"7F",x"85",x"D6",x"40",x"38",x"D3",x"FA",
x"12",x"F9",x"3C",x"FA",x"12",x"F9",x"3D",x"6F",x"E5",x"D9",x"E3",x"D5",x"C5",x"E5",
x"FD",x"E5",x"E1",x"5D",x"54",x"01",x"10",x"00",x"09",x"CD",x"E8",x"F5",x"D5",x"77",
x"2B",x"77",x"2B",x"CD",x"E8",x"F5",x"21",x"0A",x"00",x"19",x"4D",x"44",x"11",x"13",
x"00",x"19",x"D1",x"13",x"E5",x"F6",x"02",x"08",x"D9",x"0E",x"0C",x"D9",x"E1",x"E5",
x"C5",x"1A",x"D9",x"08",x"F5",x"08",x"87",x"28",x"39",x"57",x"87",x"87",x"82",x"57",
x"26",x"C0",x"1E",x"00",x"06",x"10",x"08",x"F2",x"8E",x"F5",x"1C",x"1D",x"28",x"26",
x"08",x"AF",x"18",x"0D",x"FE",x"0C",x"30",x"F8",x"08",x"D9",x"0A",x"D9",x"82",x"C6",
x"03",x"6F",x"7E",x"83",x"27",x"D9",x"86",x"27",x"36",x"00",x"ED",x"6F",x"23",x"03",
x"D9",x"07",x"07",x"07",x"07",x"5F",x"08",x"3D",x"10",x"D3",x"F1",x"3C",x"08",x"0D",
x"D9",x"C1",x"0B",x"13",x"20",x"B2",x"E1",x"01",x"0F",x"00",x"09",x"5D",x"54",x"CD",
x"DA",x"F5",x"E5",x"FD",x"E1",x"E1",x"7C",x"E6",x"80",x"B5",x"FD",x"77",x"08",x"FD",
x"36",x"00",x"09",x"C1",x"D1",x"E1",x"D9",x"C3",x"EF",x"F4",x"06",x"07",x"1A",x"1B",
x"ED",x"6F",x"1A",x"1B",x"ED",x"6F",x"2B",x"10",x"F5",x"C9",x"06",x"07",x"AF",x"ED",
x"6F",x"12",x"1B",x"AF",x"ED",x"6F",x"12",x"1B",x"2B",x"10",x"F3",x"AF",x"C9",x"CF",
x"0B",x"F5",x"FD",x"7E",x"06",x"B7",x"28",x"F7",x"FD",x"7E",x"0F",x"B7",x"CA",x"1A",
x"FA",x"D9",x"E5",x"D5",x"C5",x"FD",x"E5",x"11",x"09",x"00",x"FD",x"19",x"FD",x"6E",
x"FF",x"FD",x"66",x"08",x"E3",x"22",x"1C",x"17",x"E5",x"FD",x"E3",x"CD",x"F1",x"F9",
x"06",x"04",x"2A",x"1C",x"17",x"D9",x"01",x"F7",x"FF",x"2A",x"1C",x"17",x"5D",x"54",
x"B7",x"ED",x"42",x"EB",x"09",x"09",x"06",x"07",x"B7",x"13",x"1A",x"D9",x"23",x"9E",
x"D9",x"27",x"23",x"77",x"10",x"F5",x"E6",x"F0",x"20",x"13",x"D9",x"CD",x"D2",x"F7",
x"3C",x"CD",x"E3",x"F7",x"2A",x"1C",x"17",x"D9",x"01",x"07",x"00",x"ED",x"B8",x"18",
x"DB",x"FD",x"E3",x"CD",x"84",x"F7",x"FD",x"E3",x"D9",x"04",x"78",x"FE",x"10",x"38",
x"BB",x"D9",x"2A",x"1C",x"17",x"2B",x"2B",x"01",x"08",x"00",x"ED",x"B8",x"FD",x"E1",
x"E1",x"7C",x"AD",x"E6",x"80",x"4F",x"CB",x"BC",x"CB",x"BD",x"7C",x"95",x"C6",x"40",
x"A9",x"FD",x"77",x"08",x"A9",x"F2",x"D3",x"F5",x"CD",x"F9",x"F9",x"18",x"F8",x"FD",
x"E5",x"E1",x"01",x"09",x"00",x"09",x"5D",x"54",x"1B",x"09",x"E5",x"FD",x"E1",x"2B",
x"7E",x"E6",x"80",x"0F",x"4F",x"1A",x"E6",x"80",x"0F",x"91",x"C0",x"81",x"28",x"01",
x"EB",x"1A",x"1B",x"E6",x"7F",x"4F",x"7E",x"2B",x"E6",x"7F",x"91",x"C0",x"06",x"07",
x"1A",x"E6",x"F0",x"0F",x"4F",x"7E",x"E6",x"F0",x"0F",x"91",x"C0",x"1A",x"E6",x"0F",
x"4F",x"7E",x"E6",x"0F",x"91",x"C0",x"1B",x"2B",x"10",x"E8",x"C9",x"FD",x"E5",x"E1",
x"23",x"E5",x"4E",x"06",x"00",x"09",x"23",x"23",x"E5",x"7E",x"B9",x"38",x"01",x"79",
x"4E",x"09",x"23",x"E5",x"FD",x"E1",x"4F",x"03",x"D1",x"E1",x"1A",x"13",x"ED",x"A1",
x"E2",x"FB",x"F6",x"28",x"F7",x"2B",x"4E",x"6F",x"60",x"ED",x"42",x"7C",x"C8",x"F8",
x"3E",x"01",x"C9",x"FD",x"CB",x"08",x"7E",x"C8",x"FD",x"E5",x"E1",x"11",x"07",x"00",
x"B7",x"23",x"7A",x"9E",x"27",x"77",x"1D",x"20",x"F8",x"C9",x"FD",x"CB",x"08",x"7E",
x"C8",x"CD",x"0C",x"F7",x"18",x"05",x"FD",x"7E",x"06",x"B7",x"C8",x"3E",x"80",x"FD",
x"AE",x"08",x"FD",x"77",x"08",x"C9",x"CD",x"DF",x"F9",x"C8",x"FD",x"7E",x"07",x"B7",
x"28",x"13",x"3E",x"01",x"CD",x"90",x"F7",x"FD",x"7E",x"08",x"E6",x"7F",x"FE",x"7E",
x"CA",x"12",x"F9",x"FD",x"34",x"08",x"C9",x"FD",x"7E",x"06",x"E6",x"F0",x"C0",x"CD",
x"84",x"F7",x"FD",x"7E",x"08",x"FD",x"35",x"08",x"E6",x"7F",x"20",x"ED",x"C3",x"F9",
x"F9",x"E5",x"FD",x"E5",x"E1",x"23",x"7E",x"FE",x"50",x"36",x"00",x"38",x"0F",x"06",
x"06",x"23",x"7E",x"C6",x"01",x"27",x"77",x"30",x"02",x"10",x"F6",x"CD",x"34",x"F7",
x"E1",x"C9",x"FD",x"E5",x"E1",x"06",x"07",x"AF",x"23",x"ED",x"6F",x"10",x"FB",x"C9",
x"FE",x"0E",x"30",x"30",x"01",x"FF",x"00",x"FD",x"E5",x"E1",x"E5",x"5D",x"54",x"23",
x"D6",x"02",x"0C",x"30",x"FA",x"28",x"12",x"13",x"F5",x"3E",x"07",x"91",x"4F",x"ED",
x"B0",x"EB",x"D6",x"08",x"2F",x"70",x"23",x"3D",x"20",x"FB",x"F1",x"E1",x"3C",x"C0",
x"0E",x"07",x"09",x"41",x"ED",x"67",x"2B",x"10",x"FB",x"C9",x"FD",x"4E",x"08",x"CD",
x"F9",x"F9",x"FD",x"71",x"08",x"C9",x"21",x"B6",x"FE",x"E5",x"E5",x"C5",x"CD",x"FD",
x"F7",x"38",x"05",x"7E",x"07",x"07",x"07",x"07",x"E6",x"0F",x"C1",x"E1",x"C9",x"E5",
x"C5",x"CD",x"FD",x"F7",x"06",x"F0",x"38",x"0B",x"CB",x"21",x"CB",x"21",x"CB",x"21",
x"CB",x"21",x"7E",x"06",x"0F",x"A0",x"B1",x"77",x"C1",x"E1",x"C9",x"FD",x"E5",x"E1",
x"CB",x"38",x"F5",x"3E",x"08",x"90",x"4F",x"06",x"00",x"09",x"F1",x"4F",x"7E",x"C9",
x"FD",x"7E",x"06",x"B7",x"21",x"31",x"19",x"36",x"30",x"28",x"7E",x"FD",x"CB",x"08",
x"7E",x"28",x"06",x"36",x"2D",x"23",x"CD",x"26",x"F7",x"CD",x"67",x"F7",x"06",x"0E",
x"05",x"78",x"FE",x"04",x"D4",x"D2",x"F7",x"28",x"F7",x"48",x"06",x"04",x"FD",x"5E",
x"08",x"7B",x"D6",x"3B",x"57",x"7B",x"FE",x"4A",x"30",x"16",x"FE",x"40",x"30",x"0A",
x"91",x"38",x"10",x"FE",x"32",x"38",x"0C",x"42",x"18",x"0B",x"79",x"BA",x"30",x"07",
x"4A",x"B7",x"18",x"04",x"37",x"16",x"05",x"0C",x"F5",x"78",x"BA",x"20",x"03",x"36",
x"2E",x"23",x"78",x"D6",x"04",x"3E",x"00",x"F4",x"D2",x"F7",x"C6",x"30",x"77",x"23",
x"04",x"78",x"B9",x"20",x"E9",x"F1",x"30",x"20",x"36",x"45",x"23",x"36",x"2B",x"7B",
x"D6",x"40",x"30",x"04",x"36",x"2D",x"ED",x"44",x"23",x"06",x"FF",x"04",x"4F",x"D6",
x"0A",x"30",x"FA",x"78",x"C6",x"30",x"77",x"23",x"90",x"81",x"77",x"23",x"11",x"30",
x"19",x"37",x"ED",x"52",x"EB",x"73",x"C9",x"D5",x"C5",x"1E",x"FF",x"0E",x"00",x"7E",
x"23",x"FE",x"20",x"28",x"FA",x"FE",x"22",x"20",x"03",x"0C",x"7E",x"23",x"1C",x"0C",
x"0D",x"28",x"0E",x"FE",x"FF",x"28",x"16",x"FE",x"22",x"20",x"F1",x"BE",x"23",x"28",
x"ED",x"18",x"0C",x"FE",x"2C",x"28",x"08",x"FE",x"21",x"28",x"04",x"FE",x"FD",x"38",
x"DF",x"2B",x"E5",x"D5",x"43",x"FD",x"E5",x"D1",x"CD",x"8E",x"FC",x"04",x"05",x"1B",
x"28",x"16",x"2B",x"7E",x"FE",x"22",x"20",x"06",x"0C",x"0D",x"28",x"02",x"2B",x"7E",
x"12",x"FE",x"20",x"30",x"EB",x"F6",x"80",x"12",x"18",x"E6",x"EB",x"D1",x"73",x"2B",
x"36",x"01",x"E5",x"FD",x"E1",x"E1",x"C1",x"D1",x"C9",x"7E",x"FE",x"22",x"28",x"97",
x"CD",x"14",x"F9",x"D2",x"5A",x"FD",x"17",x"D0",x"CF",x"0D",x"C5",x"D5",x"CD",x"F4",
x"F9",x"E5",x"FD",x"E5",x"E1",x"11",x"07",x"00",x"19",x"E3",x"1E",x"3F",x"06",x"0B",
x"7E",x"23",x"FE",x"20",x"28",x"FA",x"FE",x"2B",x"28",x"06",x"FE",x"2D",x"20",x"04",
x"CB",x"CA",x"7E",x"23",x"FE",x"2E",x"28",x"2D",x"D6",x"3A",x"30",x"31",x"C6",x"0A",
x"30",x"2D",x"4F",x"CB",x"FA",x"7A",x"0F",x"20",x"09",x"CB",x"52",x"20",x"07",x"30",
x"E5",x"1D",x"18",x"E2",x"CB",x"D2",x"38",x"01",x"1C",x"78",x"3D",x"28",x"D9",x"47",
x"E3",x"0F",x"38",x"01",x"2B",x"79",x"ED",x"6F",x"E3",x"18",x"CD",x"CB",x"FA",x"CB",
x"42",x"CB",x"C2",x"28",x"C5",x"E3",x"05",x"CB",x"40",x"28",x"03",x"AF",x"ED",x"6F",
x"E1",x"2B",x"7E",x"CD",x"C8",x"FB",x"FE",x"45",x"7B",x"20",x"40",x"CB",x"FA",x"23",
x"7E",x"FE",x"98",x"28",x"0E",x"FE",x"2B",x"28",x"0A",x"FE",x"A2",x"28",x"04",x"FE",
x"2D",x"20",x"03",x"CB",x"EA",x"23",x"06",x"00",x"2B",x"23",x"7E",x"D6",x"3A",x"30",
x"12",x"C6",x"0A",x"30",x"0E",x"4F",x"78",x"87",x"47",x"87",x"87",x"80",x"81",x"47",
x"F2",x"9F",x"F9",x"CB",x"F2",x"78",x"CB",x"6A",x"28",x"02",x"ED",x"44",x"83",x"FE",
x"7F",x"38",x"02",x"CB",x"F2",x"D5",x"FD",x"77",x"08",x"CB",x"4A",x"C4",x"26",x"F7",
x"CD",x"DF",x"F9",x"D1",x"7A",x"1F",x"A2",x"E6",x"20",x"7A",x"17",x"C4",x"F9",x"F9",
x"D1",x"C1",x"C9",x"E5",x"FD",x"E5",x"E1",x"06",x"07",x"AF",x"23",x"B6",x"20",x"05",
x"10",x"FA",x"FD",x"77",x"08",x"E1",x"C9",x"CD",x"8E",x"FC",x"11",x"F7",x"FF",x"FD",
x"19",x"FD",x"E5",x"E3",x"36",x"09",x"06",x"08",x"AF",x"23",x"77",x"10",x"FC",x"E1",
x"37",x"C9",x"CD",x"F9",x"F9",x"FD",x"36",x"08",x"40",x"FD",x"36",x"06",x"10",x"C9",
x"21",x"B6",x"FE",x"E5",x"18",x"DF",x"F1",x"11",x"09",x"00",x"FD",x"19",x"C9",x"FD",
x"5E",x"01",x"16",x"00",x"13",x"13",x"FD",x"19",x"C9",x"CD",x"F1",x"F9",x"FD",x"23",
x"FD",x"22",x"1C",x"17",x"FD",x"2B",x"E5",x"CD",x"83",x"FC",x"37",x"ED",x"6A",x"30",
x"FC",x"0E",x"01",x"18",x"0F",x"04",x"0C",x"3E",x"41",x"13",x"1A",x"8F",x"27",x"12",
x"10",x"F9",x"38",x"F3",x"ED",x"6A",x"ED",x"5B",x"1C",x"17",x"20",x"EE",x"F1",x"E6",
x"80",x"F6",x"49",x"FD",x"77",x"08",x"C3",x"34",x"F7",x"CD",x"8E",x"FC",x"01",x"05",
x"00",x"09",x"FD",x"E5",x"D1",x"1B",x"ED",x"A8",x"AF",x"12",x"1B",x"03",x"ED",x"B8",
x"12",x"3E",x"09",x"1B",x"18",x"11",x"23",x"4E",x"06",x"00",x"CD",x"8E",x"FC",x"09",
x"03",x"FD",x"E5",x"D1",x"1B",x"ED",x"B8",x"3E",x"01",x"12",x"D5",x"FD",x"E1",x"C9",
x"CD",x"8E",x"FC",x"FD",x"E5",x"D1",x"1B",x"21",x"09",x"00",x"4D",x"44",x"19",x"ED",
x"B8",x"13",x"D5",x"FD",x"E1",x"C9",x"CD",x"8E",x"FC",x"FD",x"E5",x"E1",x"2B",x"5D",
x"54",x"01",x"12",x"00",x"09",x"ED",x"B8",x"13",x"D5",x"FD",x"E1",x"C9",x"CD",x"43",
x"FC",x"18",x"05",x"CD",x"C3",x"FA",x"EB",x"F6",x"37",x"C5",x"D5",x"DC",x"A7",x"F0",
x"FD",x"7E",x"08",x"F5",x"E6",x"7F",x"ED",x"62",x"FE",x"45",x"30",x"3E",x"D6",x"40",
x"38",x"2C",x"C6",x"05",x"4F",x"06",x"04",x"7C",x"E6",x"E0",x"20",x"30",x"29",x"5D",
x"54",x"29",x"29",x"19",x"38",x"28",x"CD",x"D2",x"F7",x"5F",x"16",x"00",x"19",x"38",
x"1F",x"04",x"79",x"B8",x"20",x"E5",x"F1",x"F5",x"B7",x"FC",x"86",x"FC",x"F1",x"AC",
x"FA",x"14",x"FB",x"3E",x"F1",x"11",x"09",x"00",x"FD",x"19",x"7C",x"B7",x"D9",x"78",
x"D9",x"D1",x"C1",x"C9",x"CF",x"04",x"CD",x"43",x"FC",x"3E",x"F6",x"37",x"E5",x"CD",
x"C5",x"FA",x"24",x"25",x"C2",x"14",x"FB",x"7D",x"E1",x"C9",x"CD",x"67",x"F7",x"EB",
x"FD",x"E5",x"E1",x"23",x"23",x"01",x"05",x"00",x"ED",x"B0",x"23",x"ED",x"A0",x"18",
x"1C",x"DD",x"CB",x"01",x"4E",x"20",x"E7",x"4E",x"23",x"FD",x"E5",x"D1",x"13",x"1A",
x"0C",x"20",x"01",x"0D",x"B9",x"D2",x"12",x"F9",x"4F",x"06",x"00",x"03",x"EB",x"ED",
x"B0",x"E5",x"FD",x"E1",x"C9",x"E1",x"7E",x"B7",x"E5",x"00",x"00",x"00",x"00",x"C8",
x"E1",x"C3",x"5C",x"FD",x"C3",x"00",x"00",x"C3",x"82",x"FB",x"32",x"1F",x"00",x"F7",
x"00",x"C9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"22",x"1E",x"17",x"32",x"04",x"17",x"2A",x"18",x"17",x"E3",x"7E",x"23",
x"22",x"18",x"17",x"87",x"F5",x"C6",x"C7",x"6F",x"26",x"C0",x"7E",x"23",x"66",x"6F",
x"22",x"16",x"00",x"2A",x"1E",x"17",x"3A",x"04",x"17",x"CD",x"15",x"00",x"32",x"04",
x"17",x"22",x"1E",x"17",x"2A",x"18",x"17",x"F1",x"30",x"D8",x"E3",x"22",x"18",x"17",
x"2A",x"1E",x"17",x"3A",x"04",x"17",x"C9",x"1A",x"04",x"05",x"C0",x"FE",x"FF",x"C8",
x"E6",x"7F",x"FE",x"20",x"38",x"09",x"FE",x"61",x"D8",x"FE",x"7B",x"D0",x"E6",x"DF",
x"C9",x"FE",x"10",x"D8",x"FE",x"19",x"D0",x"E6",x"EF",x"C9",x"FE",x"02",x"C2",x"5A",
x"FD",x"CD",x"C3",x"FA",x"CD",x"44",x"DD",x"D0",x"CF",x"02",x"0E",x"20",x"CD",x"FD",
x"FB",x"C0",x"FE",x"FD",x"28",x"4D",x"FE",x"FE",x"D0",x"CF",x"01",x"0E",x"20",x"DD",
x"71",x"05",x"D9",x"78",x"D9",x"FE",x"A7",x"C0",x"CD",x"16",x"FB",x"E6",x"07",x"87",
x"87",x"87",x"87",x"32",x"05",x"17",x"4F",x"AF",x"D9",x"78",x"D9",x"C9",x"DD",x"36",
x"05",x"20",x"3A",x"4E",x"0B",x"4F",x"3A",x"4D",x"0B",x"B9",x"C0",x"3C",x"32",x"4D",
x"0B",x"3A",x"13",x"0B",x"CB",x"4F",x"C8",x"79",x"2F",x"32",x"4D",x"0B",x"C9",x"DD",
x"CB",x"00",x"5E",x"C8",x"DD",x"CB",x"00",x"9E",x"F7",x"54",x"F7",x"D4",x"C9",x"D9",
x"7E",x"47",x"FE",x"FE",x"30",x"30",x"23",x"FE",x"C5",x"28",x"2F",x"FE",x"80",x"30",
x"27",x"FE",x"20",x"28",x"ED",x"2B",x"06",x"00",x"FE",x"22",x"37",x"28",x"17",x"CB",
x"C8",x"FE",x"41",x"38",x"11",x"FE",x"5B",x"3F",x"38",x"0C",x"CD",x"D2",x"F3",x"D4",
x"0B",x"F4",x"79",x"E6",x"02",x"F6",x"01",x"47",x"DC",x"05",x"F9",x"78",x"D9",x"FE",
x"FD",x"C9",x"4F",x"06",x"01",x"18",x"F6",x"CB",x"7C",x"C8",x"2B",x"7D",x"2F",x"6F",
x"7C",x"2F",x"67",x"C9",x"E5",x"D5",x"11",x"00",x"01",x"CD",x"99",x"FC",x"D1",x"E1",
x"C9",x"2A",x"26",x"17",x"19",x"38",x"12",x"EB",x"FD",x"E5",x"E1",x"ED",x"52",x"38",
x"0A",x"ED",x"62",x"39",x"ED",x"5B",x"17",x"0B",x"ED",x"52",x"D0",x"CF",x"06",x"AF",
x"6F",x"67",x"3E",x"10",x"3D",x"F8",x"ED",x"6A",x"CB",x"21",x"CB",x"10",x"30",x"F6",
x"19",x"18",x"F3",x"CD",x"D1",x"FC",x"D0",x"FE",x"CA",x"D0",x"CD",x"D5",x"FC",x"18",
x"F7",x"D9",x"E5",x"D9",x"E1",x"7E",x"FE",x"FE",x"D0",x"23",x"FE",x"FD",x"20",x"F7",
x"7E",x"23",x"FE",x"20",x"28",x"FA",x"2B",x"37",x"C9",x"06",x"00",x"FD",x"E5",x"E1",
x"4E",x"B9",x"C8",x"0C",x"0D",x"37",x"C8",x"0D",x"20",x"02",x"23",x"4E",x"0C",x"09",
x"E5",x"FD",x"E1",x"18",x"ED",x"CD",x"A7",x"F0",x"21",x"00",x"80",x"E5",x"CD",x"2B",
x"FA",x"CD",x"93",x"F4",x"CD",x"C3",x"FA",x"D1",x"19",x"C9",x"4F",x"7E",x"B7",x"79",
x"C8",x"96",x"23",x"5E",x"23",x"20",x"F6",x"57",x"19",x"CD",x"43",x"FC",x"CD",x"AD",
x"DB",x"37",x"C9",x"CD",x"43",x"FC",x"1E",x"01",x"28",x"08",x"CD",x"45",x"FD",x"5A",
x"FE",x"FD",x"20",x"0A",x"CD",x"43",x"FC",x"16",x"FF",x"FE",x"95",x"C4",x"45",x"FD",
x"3E",x"95",x"C3",x"54",x"FD",x"CD",x"C4",x"FA",x"16",x"00",x"24",x"C8",x"15",x"25",
x"C0",x"55",x"C9",x"CD",x"43",x"FC",x"D9",x"B8",x"D9",x"CA",x"43",x"FC",x"3E",x"01",
x"FD",x"2A",x"1A",x"17",x"FE",x"F5",x"CA",x"A3",x"FF",x"F5",x"FE",x"06",x"CC",x"FC",
x"DC",x"CD",x"35",x"FC",x"CD",x"18",x"FC",x"CD",x"79",x"FE",x"06",x"0D",x"0A",x"2A",
x"2A",x"2A",x"20",x"F1",x"CB",x"7F",x"20",x"18",x"21",x"C6",x"FD",x"01",x"FF",x"FF",
x"03",x"09",x"4E",x"23",x"0C",x"0D",x"28",x"04",x"B9",x"4E",x"20",x"F4",x"23",x"CD",
x"DD",x"FE",x"18",x"18",x"6F",x"CD",x"79",x"FE",x"0D",x"53",x"79",x"73",x"74",x"65",
x"6D",x"20",x"65",x"72",x"72",x"6F",x"72",x"20",x"AF",x"67",x"47",x"CD",x"1B",x"FF",
x"CD",x"79",x"FE",x"04",x"2E",x"0B",x"0D",x"0A",x"DD",x"CB",x"00",x"CE",x"2A",x"0C",
x"17",x"AF",x"CD",x"2D",x"DD",x"C3",x"0E",x"E1",x"01",x"0F",x"4E",x"6F",x"74",x"20",
x"75",x"6E",x"64",x"65",x"72",x"73",x"74",x"6F",x"6F",x"64",x"FF",x"02",x"06",x"4C",
x"69",x"6E",x"65",x"93",x"FF",x"03",x"04",x"41",x"92",x"93",x"FF",x"04",x"04",x"91",
x"61",x"92",x"FF",x"05",x"0B",x"91",x"73",x"75",x"62",x"73",x"63",x"72",x"69",x"70",
x"74",x"FF",x"06",x"08",x"90",x"6D",x"65",x"6D",x"6F",x"72",x"79",x"FF",x"07",x"03",
x"90",x"FB",x"FF",x"08",x"03",x"90",x"F2",x"FF",x"09",x"03",x"90",x"F0",x"FF",x"0A",
x"03",x"8F",x"F8",x"FF",x"0B",x"0D",x"8F",x"64",x"69",x"76",x"69",x"64",x"65",x"20",
x"62",x"79",x"20",x"30",x"FF",x"0C",x"03",x"8F",x"DB",x"FF",x"0D",x"09",x"4F",x"76",
x"65",x"72",x"66",x"6C",x"6F",x"77",x"FF",x"0E",x"0E",x"54",x"79",x"70",x"65",x"20",
x"6D",x"69",x"73",x"6D",x"61",x"74",x"63",x"68",x"FF",x"0F",x"18",x"56",x"61",x"72",
x"69",x"61",x"62",x"6C",x"65",x"20",x"64",x"65",x"63",x"6C",x"61",x"72",x"65",x"64",
x"20",x"74",x"77",x"69",x"63",x"65",x"FF",x"10",x"06",x"91",x"66",x"69",x"6C",x"65",
x"FF",x"00",x"0F",x"42",x"41",x"53",x"49",x"43",x"20",x"63",x"6F",x"72",x"72",x"75",
x"70",x"74",x"65",x"64",x"FF",x"E3",x"CD",x"7F",x"FE",x"E3",x"C9",x"7E",x"23",x"B7",
x"C8",x"C5",x"47",x"7E",x"23",x"CD",x"9A",x"FE",x"10",x"F9",x"C1",x"C9",x"3E",x"0B",
x"CC",x"9A",x"FE",x"3E",x"0D",x"CD",x"9A",x"FE",x"3E",x"0A",x"F5",x"C5",x"D5",x"4F",
x"CD",x"A6",x"FE",x"D7",x"D1",x"C1",x"F1",x"C9",x"11",x"7F",x"00",x"3A",x"05",x"17",
x"F6",x"01",x"B2",x"A3",x"C3",x"1B",x"00",x"CD",x"9A",x"FE",x"E1",x"C3",x"F0",x"FF",
x"FD",x"CB",x"08",x"7E",x"CC",x"C7",x"FE",x"CD",x"0E",x"F8",x"CD",x"7F",x"FE",x"3E",
x"20",x"18",x"CF",x"87",x"FE",x"40",x"1F",x"CD",x"9A",x"FE",x"FE",x"22",x"20",x"09",
x"B9",x"28",x"02",x"41",x"0E",x"78",x"0E",x"AF",x"4F",x"7E",x"23",x"3C",x"C8",x"3D",
x"F2",x"CB",x"FE",x"E5",x"0C",x"0D",x"F5",x"FE",x"FB",x"28",x"04",x"FE",x"FC",x"38",
x"02",x"0E",x"FF",x"FE",x"FD",x"20",x"03",x"F1",x"0C",x"F5",x"F1",x"20",x"12",x"2F",
x"21",x"6D",x"DE",x"CB",x"7E",x"23",x"28",x"FB",x"3D",x"20",x"F8",x"7E",x"23",x"CB",
x"7F",x"CB",x"BF",x"CD",x"9A",x"FE",x"28",x"F5",x"E1",x"18",x"C6",x"06",x"FF",x"9F",
x"E6",x"20",x"4F",x"E5",x"21",x"47",x"FF",x"5E",x"23",x"56",x"23",x"E3",x"AF",x"ED",
x"52",x"3C",x"30",x"FB",x"19",x"3D",x"28",x"07",x"0E",x"30",x"81",x"CD",x"9A",x"FE",
x"79",x"A9",x"C4",x"9A",x"FE",x"E3",x"1D",x"20",x"E2",x"E1",x"79",x"A0",x"20",x"81",
x"C9",x"E8",x"03",x"64",x"00",x"0A",x"00",x"01",x"00",x"21",x"31",x"18",x"E5",x"06",
x"00",x"C5",x"11",x"FF",x"80",x"CD",x"A9",x"FE",x"D1",x"42",x"28",x"12",x"E1",x"06",
x"00",x"70",x"23",x"36",x"FF",x"2B",x"FE",x"F5",x"28",x"2F",x"FE",x"EC",x"28",x"2B",
x"B7",x"D7",x"3A",x"16",x"0B",x"B7",x"3E",x"F5",x"20",x"E6",x"79",x"FE",x"0D",x"28",
x"13",x"FE",x"20",x"38",x"D2",x"D6",x"80",x"38",x"05",x"FE",x"20",x"30",x"01",x"4F",
x"78",x"FE",x"FB",x"30",x"C4",x"04",x"23",x"71",x"20",x"BF",x"36",x"FF",x"AF",x"E1",
x"70",x"B7",x"C9",x"3A",x"16",x"0B",x"B7",x"C8",x"D9",x"D9",x"AF",x"32",x"16",x"0B",
x"CD",x"35",x"FC",x"CD",x"18",x"FC",x"CD",x"79",x"FE",x"06",x"0D",x"0A",x"53",x"54",
x"4F",x"50",x"DD",x"CB",x"00",x"56",x"28",x"22",x"22",x"10",x"17",x"2A",x"0C",x"17",
x"22",x"0E",x"17",x"CD",x"79",x"FE",x"09",x"20",x"61",x"74",x"20",x"6C",x"69",x"6E",
x"65",x"20",x"2A",x"0C",x"17",x"23",x"5E",x"23",x"56",x"EB",x"B7",x"CD",x"19",x"FF",
x"AF",x"CD",x"8E",x"FE",x"C3",x"DA",x"DA",x"7C",x"FE",x"C0",x"D8",x"CB",x"B4",x"3E",
x"50",x"C9",x"F5",x"3E",x"F0",x"32",x"03",x"00",x"D3",x"02",x"F1",x"E9",x"79",x"FE",
x"0D",x"28",x"13",x"FE"

  );

signal  do : std_logic_vector(7 downto 0);

begin

  process(CLK)
  begin
    if rising_edge(CLK) then
	   do <= myROM(conv_integer(A));
	 end if;
  end process;  
  DOUT <= do;
  
end Behavioral;
